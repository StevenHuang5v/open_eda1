VERSION	5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
    DATABASE MICRONS 2000 ;
END UNITS

LAYER TEXT
    TYPE MASTERSLICE ;
END TEXT

LAYER PO
    TYPE MASTERSLICE ;
END PO

LAYER CO
    TYPE CUT ;
END CO

LAYER M1
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    PITCH 0.200 ;
    WIDTH 0.09 ;
    MINWIDTH 0.09 ;
    SPACING 0.09 ;
    AREA 0.042 ;
END M1

LAYER VIA1
    TYPE CUT ;
    SPACING 0.10 ;
END VIA1

LAYER M2
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    PITCH 0.200 ;
    WIDTH 0.1 ;
    MINWIDTH 0.1 ;
    SPACING 0.10 ;
    AREA 0.052 ;
END M2

LAYER VIA2
    TYPE CUT ;
    SPACING 0.10 ;
END VIA2

LAYER M3
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    PITCH 0.200 ;
    WIDTH 0.1 ;
    MINWIDTH 0.1 ;
    SPACING 0.10 ;
    AREA 0.052 ;
END M3

LAYER VIA3
    TYPE CUT ;
    SPACING 0.10 ;
END VIA3

LAYER M4
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    PITCH 0.200 ;
    WIDTH 0.1 ;
    MINWIDTH 0.1 ;
    SPACING 0.10 ;
    AREA 0.052 ;
END M4

LAYER VIA4
    TYPE CUT ;
    SPACING 0.10 ;
END VIA4

LAYER M5
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    PITCH 0.200 ;
    WIDTH 0.1 ;
    MINWIDTH 0.1 ;
    SPACING 0.10 ;
    AREA 0.052 ;
END M5

LAYER VIA5
    TYPE CUT ;
    SPACING 0.340 ;
END VIA5

LAYER M6
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    PITCH 0.800 ;
    WIDTH 0.400 ;
    MINWIDTH 0.400 ;
    SPACING 0.40 ;
    AREA 0.565 ;
END M6

VIA VIA12_1cut DEFAULT
    LAYER M1 ;
        RECT -0.090 -0.050  0.090  0.050 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M2 ;
        RECT -0.050 -0.090  0.050  0.090 ;
END VIA12_1cut

VIA VIA12_1cut_H DEFAULT
    LAYER M1 ;
        RECT -0.090 -0.050  0.090  0.050 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M2 ;
        RECT -0.090 -0.050  0.090  0.050 ;
END VIA12_1cut_H
                 
VIA VIA12_1cut_V DEFAULT
    LAYER M1 ;
        RECT -0.050 -0.090  0.050  0.090 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M2 ;
        RECT -0.050 -0.090  0.050  0.090 ;
END VIA12_1cut_V

VIA VIA12_1cut_FAT_C DEFAULT
    LAYER M1 ;
        RECT -0.12 -0.050  0.12  0.050 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M2 ;
        RECT -0.050 -0.12  0.050  0.12 ;
END VIA12_1cut_FAT_C
             
VIA VIA12_1cut_FAT_H DEFAULT
    LAYER M1 ;
        RECT -0.12 -0.050  0.12  0.050 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M2 ;
        RECT -0.12 -0.050  0.12  0.050 ;
END VIA12_1cut_FAT_H

VIA VIA12_1cut_FAT_V DEFAULT
    LAYER M1 ;
        RECT -0.050 -0.12  0.050  0.12 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M2 ;
        RECT -0.050 -0.12  0.050  0.12 ;
END VIA12_1cut_FAT_V

VIA VIA12_1cut_FAT DEFAULT
    LAYER M1 ;
        RECT -0.080 -0.080  0.080  0.080 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M2 ;
        RECT -0.080 -0.080  0.080  0.080 ;
END VIA12_1cut_FAT
                 
VIA VIA12_2cut_E DEFAULT
    LAYER M1 ;
        RECT -0.090 -0.050  0.290  0.050 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT  0.150 -0.050  0.250  0.050 ;
    LAYER M2 ;
        RECT -0.050 -0.090  0.250  0.090 ;
END VIA12_2cut_E

VIA VIA12_2cut_W DEFAULT
    LAYER M1 ;
        RECT -0.290 -0.050  0.090  0.050 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.250 -0.050 -0.150  0.050 ;
    LAYER M2 ;
        RECT -0.250 -0.090  0.050  0.090 ;
END VIA12_2cut_W

VIA VIA12_2cut_N DEFAULT
    LAYER M1 ;
        RECT -0.090 -0.050  0.090  0.250 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050  0.150  0.050  0.250 ;
    LAYER M2 ;
        RECT -0.050 -0.090  0.050  0.290 ;
END VIA12_2cut_N

VIA VIA12_2cut_S DEFAULT
    LAYER M1 ;
        RECT -0.090 -0.250  0.090  0.050 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050 -0.250  0.050 -0.150 ;
    LAYER M2 ;
        RECT -0.050 -0.290  0.050  0.090 ;
END VIA12_2cut_S

VIA VIA12_2cut_HN DEFAULT
    LAYER M1 ;
        RECT -0.050 -0.090  0.050  0.330 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050  0.190  0.050  0.290 ;
    LAYER M2 ;
        RECT -0.050 -0.090  0.050  0.330 ;
END VIA12_2cut_HN

VIA VIA12_2cut_HS DEFAULT
    LAYER M1 ;
        RECT -0.050 -0.330  0.050  0.090 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050 -0.290  0.050 -0.190 ;
    LAYER M2 ;
        RECT -0.050 -0.330  0.050  0.090 ;
END VIA12_2cut_HS

VIA VIA12_4cut DEFAULT
    LAYER M1 ;
        RECT -0.190 -0.150  0.190  0.150 ;
    LAYER VIA1 ;
        RECT -0.150 -0.150 -0.050 -0.050 ;
        RECT -0.150  0.050 -0.050  0.150 ;
        RECT  0.050  0.050  0.150  0.150 ;
        RECT  0.050 -0.150  0.150 -0.050 ;
    LAYER M2 ;
        RECT -0.150 -0.190  0.150  0.190 ;
END VIA12_4cut

VIA VIA23_1cut DEFAULT
    LAYER M2 ;
        RECT -0.050 -0.090  0.050  0.090 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M3 ;
        RECT -0.090 -0.050  0.090  0.050 ;
END VIA23_1cut

VIA VIA23_1cut_V DEFAULT
    LAYER M2 ;
        RECT -0.050 -0.090  0.050  0.090 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M3 ;
        RECT -0.050 -0.090  0.050  0.090 ;
END VIA23_1cut_V
                 
VIA VIA23_1cut_H DEFAULT
    LAYER M2 ;
        RECT -0.090 -0.050  0.090  0.050 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M3 ;
        RECT -0.090 -0.050  0.090  0.050 ;
END VIA23_1cut_H

VIA VIA23_1cut_FAT_C DEFAULT
    LAYER M2 ;
        RECT -0.050 -0.12  0.050  0.12 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M3 ;
        RECT -0.12 -0.050  0.12  0.050 ;
END VIA23_1cut_FAT_C
             
VIA VIA23_1cut_FAT_V DEFAULT
    LAYER M2 ;
        RECT -0.050 -0.12  0.050  0.12 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M3 ;
        RECT -0.050 -0.12  0.050  0.12 ;
END VIA23_1cut_FAT_V

VIA VIA23_1cut_FAT_H DEFAULT
    LAYER M2 ;
        RECT -0.12 -0.050  0.12  0.050 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M3 ;
        RECT -0.12 -0.050  0.12  0.050 ;
END VIA23_1cut_FAT_H

VIA VIA23_1cut_FAT DEFAULT
    LAYER M2 ;
        RECT -0.080 -0.080  0.080  0.080 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M3 ;
        RECT -0.080 -0.080  0.080  0.080 ;
END VIA23_1cut_FAT
                 
VIA VIA23_1stack_N DEFAULT
    LAYER M2 ;
        RECT -0.050 -0.090  0.050  0.430 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M3 ;
        RECT -0.090 -0.050  0.090  0.050 ;
END VIA23_1stack_N

VIA VIA23_1stack_S DEFAULT
    LAYER M2 ;
        RECT -0.050 -0.430  0.050  0.090 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M3 ;
        RECT -0.090 -0.050  0.090  0.050 ;
END VIA23_1stack_S

VIA VIA23_2cut_E DEFAULT
    LAYER M2 ;
        RECT -0.050 -0.090  0.250  0.090 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT  0.150 -0.050  0.250  0.050 ;
    LAYER M3 ;
        RECT -0.090 -0.050  0.290  0.050 ;
END VIA23_2cut_E

VIA VIA23_2cut_W DEFAULT
    LAYER M2 ;
        RECT -0.250 -0.090  0.050  0.090 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.250 -0.050 -0.150  0.050 ;
    LAYER M3 ;
        RECT -0.290 -0.050  0.090  0.050 ;
END VIA23_2cut_W

VIA VIA23_2cut_N DEFAULT
    LAYER M2 ;
        RECT -0.050 -0.090  0.050  0.290 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050  0.150  0.050  0.250 ;
    LAYER M3 ;
        RECT -0.090 -0.050  0.090  0.250 ;
END VIA23_2cut_N

VIA VIA23_2cut_S DEFAULT
    LAYER M2 ;
        RECT -0.050 -0.290  0.050  0.090 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050 -0.250  0.050 -0.150 ;
    LAYER M3 ;
        RECT -0.090 -0.250  0.090  0.050 ;
END VIA23_2cut_S

VIA VIA23_4cut DEFAULT
    LAYER M2 ;
        RECT -0.150 -0.190  0.150  0.190 ;
    LAYER VIA2 ;
        RECT -0.150 -0.150 -0.050 -0.050 ;
        RECT -0.150  0.050 -0.050  0.150 ;
        RECT  0.050  0.050  0.150  0.150 ;
        RECT  0.050 -0.150  0.150 -0.050 ;
    LAYER M3 ;
        RECT -0.190 -0.150  0.190  0.150 ;
END VIA23_4cut

VIA VIA34_1cut DEFAULT
    LAYER M3 ;
        RECT -0.090 -0.050  0.090  0.050 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M4 ;
        RECT -0.050 -0.090  0.050  0.090 ;
END VIA34_1cut

VIA VIA34_1cut_H DEFAULT
    LAYER M3 ;
        RECT -0.090 -0.050  0.090  0.050 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M4 ;
        RECT -0.090 -0.050  0.090  0.050 ;
END VIA34_1cut_H
                 
VIA VIA34_1cut_V DEFAULT
    LAYER M3 ;
        RECT -0.050 -0.090  0.050  0.090 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M4 ;
        RECT -0.050 -0.090  0.050  0.090 ;
END VIA34_1cut_V

VIA VIA34_1cut_FAT_C DEFAULT
    LAYER M3 ;
        RECT -0.12 -0.050  0.12  0.050 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M4 ;
        RECT -0.050 -0.12  0.050  0.12 ;
END VIA34_1cut_FAT_C
             
VIA VIA34_1cut_FAT_H DEFAULT
    LAYER M3 ;
        RECT -0.12 -0.050  0.12  0.050 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M4 ;
        RECT -0.12 -0.050  0.12  0.050 ;
END VIA34_1cut_FAT_H

VIA VIA34_1cut_FAT_V DEFAULT
    LAYER M3 ;
        RECT -0.050 -0.12  0.050  0.12 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M4 ;
        RECT -0.050 -0.12  0.050  0.12 ;
END VIA34_1cut_FAT_V

VIA VIA34_1cut_FAT DEFAULT
    LAYER M3 ;
        RECT -0.080 -0.080  0.080  0.080 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M4 ;
        RECT -0.080 -0.080  0.080  0.080 ;
END VIA34_1cut_FAT
                 
VIA VIA34_1stack_E DEFAULT
    LAYER M3 ;
        RECT -0.090 -0.050  0.430  0.050 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M4 ;
        RECT -0.050 -0.090  0.050  0.090 ;
END VIA34_1stack_E

VIA VIA34_1stack_W DEFAULT
    LAYER M3 ;
        RECT -0.430 -0.050  0.090  0.050 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M4 ;
        RECT -0.050 -0.090  0.050  0.090 ;
END VIA34_1stack_W

VIA VIA34_2cut_E DEFAULT
    LAYER M3 ;
        RECT -0.090 -0.050  0.290  0.050 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT  0.150 -0.050  0.250  0.050 ;
    LAYER M4 ;
        RECT -0.050 -0.090  0.250  0.090 ;
END VIA34_2cut_E

VIA VIA34_2cut_W DEFAULT
    LAYER M3 ;
        RECT -0.290 -0.050  0.090  0.050 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.250 -0.050 -0.150  0.050 ;
    LAYER M4 ;
        RECT -0.250 -0.090  0.050  0.090 ;
END VIA34_2cut_W

VIA VIA34_2cut_N DEFAULT
    LAYER M3 ;
        RECT -0.090 -0.050  0.090  0.250 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050  0.150  0.050  0.250 ;
    LAYER M4 ;
        RECT -0.050 -0.090  0.050  0.290 ;
END VIA34_2cut_N

VIA VIA34_2cut_S DEFAULT
    LAYER M3 ;
        RECT -0.090 -0.250  0.090  0.050 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050 -0.250  0.050 -0.150 ;
    LAYER M4 ;
        RECT -0.050 -0.290  0.050  0.090 ;
END VIA34_2cut_S

VIA VIA34_4cut DEFAULT
    LAYER M3 ;
        RECT -0.190 -0.150  0.190  0.150 ;
    LAYER VIA3 ;
        RECT -0.150 -0.150 -0.050 -0.050 ;
        RECT -0.150  0.050 -0.050  0.150 ;
        RECT  0.050  0.050  0.150  0.150 ;
        RECT  0.050 -0.150  0.150 -0.050 ;
    LAYER M4 ;
        RECT -0.150 -0.190  0.150  0.190 ;
END VIA34_4cut

VIA VIA45_1cut DEFAULT
    LAYER M4 ;
        RECT -0.050 -0.090  0.050  0.090 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M5 ;
        RECT -0.090 -0.050  0.090  0.050 ;
END VIA45_1cut

VIA VIA45_1cut_V DEFAULT
    LAYER M4 ;
        RECT -0.050 -0.090  0.050  0.090 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M5 ;
        RECT -0.050 -0.090  0.050  0.090 ;
END VIA45_1cut_V
                 
VIA VIA45_1cut_H DEFAULT
    LAYER M4 ;
        RECT -0.090 -0.050  0.090  0.050 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M5 ;
        RECT -0.090 -0.050  0.090  0.050 ;
END VIA45_1cut_H

VIA VIA45_1cut_FAT_C DEFAULT
    LAYER M4 ;
        RECT -0.050 -0.12  0.050  0.12 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M5 ;
        RECT -0.12 -0.050  0.12  0.050 ;
END VIA45_1cut_FAT_C
             
VIA VIA45_1cut_FAT_V DEFAULT
    LAYER M4 ;
        RECT -0.050 -0.12  0.050  0.12 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M5 ;
        RECT -0.050 -0.12  0.050  0.12 ;
END VIA45_1cut_FAT_V

VIA VIA45_1cut_FAT_H DEFAULT
    LAYER M4 ;
        RECT -0.12 -0.050  0.12  0.050 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M5 ;
        RECT -0.12 -0.050  0.12  0.050 ;
END VIA45_1cut_FAT_H

VIA VIA45_1cut_FAT DEFAULT
    LAYER M4 ;
        RECT -0.080 -0.080  0.080  0.080 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M5 ;
        RECT -0.080 -0.080  0.080  0.080 ;
END VIA45_1cut_FAT
                 
VIA VIA45_1stack_N DEFAULT
    LAYER M4 ;
        RECT -0.050 -0.090  0.050  0.430 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M5 ;
        RECT -0.090 -0.050  0.090  0.050 ;
END VIA45_1stack_N

VIA VIA45_1stack_S DEFAULT
    LAYER M4 ;
        RECT -0.050 -0.430  0.050  0.090 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M5 ;
        RECT -0.090 -0.050  0.090  0.050 ;
END VIA45_1stack_S

VIA VIA45_2cut_E DEFAULT
    LAYER M4 ;
        RECT -0.050 -0.090  0.250  0.090 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT  0.150 -0.050  0.250  0.050 ;
    LAYER M5 ;
        RECT -0.090 -0.050  0.290  0.050 ;
END VIA45_2cut_E

VIA VIA45_2cut_W DEFAULT
    LAYER M4 ;
        RECT -0.250 -0.090  0.050  0.090 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.250 -0.050 -0.150  0.050 ;
    LAYER M5 ;
        RECT -0.290 -0.050  0.090  0.050 ;
END VIA45_2cut_W

VIA VIA45_2cut_N DEFAULT
    LAYER M4 ;
        RECT -0.050 -0.090  0.050  0.290 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050  0.150  0.050  0.250 ;
    LAYER M5 ;
        RECT -0.090 -0.050  0.090  0.250 ;
END VIA45_2cut_N

VIA VIA45_2cut_S DEFAULT
    LAYER M4 ;
        RECT -0.050 -0.290  0.050  0.090 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050 -0.250  0.050 -0.150 ;
    LAYER M5 ;
        RECT -0.090 -0.250  0.090  0.050 ;
END VIA45_2cut_S

VIA VIA45_2stack_N DEFAULT
    LAYER M4 ;
        RECT -0.050 -0.090  0.050  0.430 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050  0.150  0.050  0.250 ;
    LAYER M5 ;
        RECT -0.090 -0.050  0.090  0.250 ;
END VIA45_2stack_N
 
VIA VIA45_2stack_S DEFAULT
    LAYER M4 ;
        RECT -0.050 -0.430  0.050  0.090 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050 -0.250  0.050 -0.150 ;
    LAYER M5 ;
        RECT -0.090 -0.250  0.090  0.050 ;
END VIA45_2stack_S

VIA VIA45_4cut DEFAULT
    LAYER M4 ;
        RECT -0.150 -0.190  0.150  0.190 ;
    LAYER VIA4 ;
        RECT -0.150 -0.150 -0.050 -0.050 ;
        RECT -0.150  0.050 -0.050  0.150 ;
        RECT  0.050  0.050  0.150  0.150 ;
        RECT  0.050 -0.150  0.150 -0.050 ;
    LAYER M5 ;
        RECT -0.190 -0.150  0.190  0.150 ;
END VIA45_4cut

VIA VIA56_1cut DEFAULT
    LAYER M5 ;
        RECT -0.260 -0.200  0.260  0.200 ;
    LAYER VIA5 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M6 ;
        RECT -0.200 -0.260  0.200  0.260 ;
END VIA56_1cut

VIA VIA56_1cut_H DEFAULT
    LAYER M5 ;
        RECT -0.260 -0.200  0.260  0.200 ;
    LAYER VIA5 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M6 ;
        RECT -0.260 -0.200  0.260  0.200 ;
END VIA56_1cut_H
                 
VIA VIA56_1cut_V DEFAULT
    LAYER M5 ;
        RECT -0.200 -0.260  0.200  0.260 ;
    LAYER VIA5 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M6 ;
        RECT -0.200 -0.260  0.200  0.260 ;
END VIA56_1cut_V

VIA VIA56_1cut_FAT_C DEFAULT
    LAYER M5 ;
        RECT -0.26 -0.200  0.26  0.200 ;
    LAYER VIA5 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M6 ;
        RECT -0.200 -0.26  0.200  0.26 ;
END VIA56_1cut_FAT_C
             
VIA VIA56_1cut_FAT_H DEFAULT
    LAYER M5 ;
        RECT -0.26 -0.200  0.26  0.200 ;
    LAYER VIA5 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M6 ;
        RECT -0.26 -0.200  0.26  0.200 ;
END VIA56_1cut_FAT_H

VIA VIA56_1cut_FAT_V DEFAULT
    LAYER M5 ;
        RECT -0.200 -0.26  0.200  0.26 ;
    LAYER VIA5 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M6 ;
        RECT -0.200 -0.26  0.200  0.26 ;
END VIA56_1cut_FAT_V

VIA VIA56_1cut_FAT DEFAULT
    LAYER M5 ;
        RECT -0.260 -0.260  0.260  0.260 ;
    LAYER VIA5 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M6 ;
        RECT -0.260 -0.260  0.260  0.260 ;
END VIA56_1cut_FAT
                 
VIA VIA56_2cut_E DEFAULT
    LAYER M5 ;
        RECT -0.260 -0.200  0.960  0.200 ;
    LAYER VIA5 ;
        RECT -0.180 -0.180  0.180  0.180 ;
        RECT  0.520 -0.180  0.880  0.180 ;
    LAYER M6 ;
        RECT -0.200 -0.260  0.900  0.260 ;
END VIA56_2cut_E

VIA VIA56_2cut_W DEFAULT
    LAYER M5 ;
        RECT -0.960 -0.200  0.260  0.200 ;
    LAYER VIA5 ;
        RECT -0.180 -0.180  0.180  0.180 ;
        RECT -0.880 -0.180 -0.520  0.180 ;
    LAYER M6 ;
        RECT -0.900 -0.260  0.200  0.260 ;
END VIA56_2cut_W

VIA VIA56_2cut_N DEFAULT
    LAYER M5 ;
        RECT -0.260 -0.200  0.260  0.900 ;
    LAYER VIA5 ;
        RECT -0.180 -0.180  0.180  0.180 ;
        RECT -0.180  0.520  0.180  0.880 ;
    LAYER M6 ;
        RECT -0.200 -0.260  0.200  0.960 ;
END VIA56_2cut_N

VIA VIA56_2cut_S DEFAULT
    LAYER M5 ;
        RECT -0.260 -0.900  0.260  0.200 ;
    LAYER VIA5 ;
        RECT -0.180 -0.180  0.180  0.180 ;
        RECT -0.180 -0.880  0.180 -0.520 ;
    LAYER M6 ;
        RECT -0.200 -0.960  0.200  0.260 ;
END VIA56_2cut_S

VIA VIA56_4cut DEFAULT
    LAYER M5 ;
        RECT -0.710 -0.650  0.710  0.650 ;
    LAYER VIA5 ;
        RECT -0.630 -0.630 -0.270 -0.270 ;
        RECT -0.630  0.270 -0.270  0.630 ;
        RECT  0.270  0.270  0.630  0.630 ;
        RECT  0.270 -0.630  0.630 -0.270 ;
    LAYER M6 ;
        RECT -0.650 -0.710  0.650  0.710 ;
END VIA56_4cut

VIARULE VIAGEN12 GENERATE
    LAYER M1 ;
        ENCLOSURE 0.4E-01 0 ; 
        WIDTH 0.09 TO 12.00 ;
    LAYER M2 ;
        ENCLOSURE 0.4E-01 0 ;
        WIDTH 0.10 TO 12.00 ;
    LAYER VIA1 ;
        RECT -0.5E-01 -0.5E-01 0.5E-01 0.5E-01 ;
        SPACING 0.23 BY 0.23 ;    
END VIAGEN12        

VIARULE VIAGEN23 GENERATE
    LAYER M2 ;
        ENCLOSURE 0.4E-01 0 ;  
        WIDTH 0.10 TO 12.00 ;
    LAYER M3 ;
        ENCLOSURE 0.4E-01 0 ; 
        WIDTH 0.10 TO 12.00 ;
    LAYER VIA2 ;
        RECT -0.5E-01 -0.5E-01 0.5E-01 0.5E-01 ; 
        SPACING 0.23 BY 0.23 ;    
END VIAGEN23

VIARULE VIAGEN34 GENERATE
    LAYER M3 ;
        ENCLOSURE 0.4E-01 0 ; 
        WIDTH 0.10 TO 12.00 ;
    LAYER M4 ;
        ENCLOSURE 0.4E-01 0 ; 
        WIDTH 0.10 TO 12.00 ;
    LAYER VIA3 ;
        RECT -0.5E-01 -0.5E-01 0.5E-01 0.5E-01 ; 
        SPACING 0.23 BY 0.23 ;    
END VIAGEN34

VIARULE VIAGEN45 GENERATE
    LAYER M4 ;
        ENCLOSURE 0.4E-01 0 ; 
        WIDTH 0.10 TO 12.00 ;
    LAYER M5 ;
        ENCLOSURE 0.4E-01 0 ; 
        WIDTH 0.10 TO 12.00 ;
    LAYER VIA4 ;
        RECT -0.5E-01 -0.5E-01 0.5E-01 0.5E-01 ; 
        SPACING 0.23 BY 0.23 ;    
END VIAGEN45

VIARULE VIAGEN56 GENERATE
    LAYER M5 ;
        ENCLOSURE 0.8E-01 0.2E-01  ;
        WIDTH 0.10 TO 12.00 ;
    LAYER M6 ;
        ENCLOSURE 0.8E-01 0.2E-01  ;
        WIDTH 0.40 TO 12.00 ;
    LAYER VIA5 ;
        RECT -0.18 -0.18 0.18 0.18 ; 
        SPACING 0.90 BY 0.90 ;    
END VIAGEN56

MACRO CELL47
    CLASS CORE ;
    FOREIGN CELL47 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 0.1512 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.510 1.150 1.800 ;
        RECT  0.980 0.510 1.050 0.690 ;
        RECT  0.980 1.400 1.050 1.800 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0507 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 1.000 0.640 1.170 ;
        RECT  0.450 1.000 0.550 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.910 0.355 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.795 -0.330 1.200 0.330 ;
        RECT  0.645 -0.330 0.795 0.480 ;
        RECT  0.000 -0.330 0.645 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.800 2.070 1.200 2.730 ;
        RECT  0.690 1.600 0.800 2.730 ;
        RECT  0.220 2.070 0.690 2.730 ;
        RECT  0.110 1.400 0.220 2.730 ;
        RECT  0.000 2.070 0.110 2.730 ;
        END
    END VDD
END CELL47

MACRO CELL24
    CLASS CORE ;
    FOREIGN CELL24 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 0.6720 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.950 0.510 2.060 0.890 ;
        RECT  1.950 1.305 2.060 1.890 ;
        RECT  1.850 0.710 1.950 0.890 ;
        RECT  1.850 1.305 1.950 1.490 ;
        RECT  1.550 0.710 1.850 1.490 ;
        RECT  1.500 0.710 1.550 0.890 ;
        RECT  1.500 1.305 1.550 1.490 ;
        RECT  1.390 0.510 1.500 0.890 ;
        RECT  1.390 1.305 1.500 1.890 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.2018 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.985 0.960 1.100 1.180 ;
        RECT  0.750 0.960 0.985 1.070 ;
        RECT  0.650 0.690 0.750 1.070 ;
        RECT  0.360 0.690 0.650 0.780 ;
        RECT  0.270 0.690 0.360 1.000 ;
        RECT  0.180 0.910 0.270 1.000 ;
        RECT  0.050 0.910 0.180 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2019 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.890 0.550 1.310 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.325 -0.330 2.400 0.330 ;
        RECT  2.215 -0.330 2.325 0.800 ;
        RECT  1.780 -0.330 2.215 0.330 ;
        RECT  1.670 -0.330 1.780 0.600 ;
        RECT  1.230 -0.330 1.670 0.330 ;
        RECT  1.120 -0.330 1.230 0.600 ;
        RECT  0.180 -0.330 1.120 0.330 ;
        RECT  0.070 -0.330 0.180 0.800 ;
        RECT  0.000 -0.330 0.070 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.325 2.070 2.400 2.730 ;
        RECT  2.215 1.400 2.325 2.730 ;
        RECT  1.780 2.070 2.215 2.730 ;
        RECT  1.670 1.600 1.780 2.730 ;
        RECT  1.230 2.070 1.670 2.730 ;
        RECT  1.120 1.620 1.230 2.730 ;
        RECT  0.710 2.070 1.120 2.730 ;
        RECT  0.600 1.620 0.710 2.730 ;
        RECT  0.190 2.070 0.600 2.730 ;
        RECT  0.080 1.400 0.190 2.730 ;
        RECT  0.000 2.070 0.080 2.730 ;
        END
    END VDD
END CELL24

MACRO CELL91
    CLASS CORE ;
    FOREIGN CELL91 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 0.2880 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.510 1.150 1.890 ;
        RECT  0.980 0.510 1.050 0.890 ;
        RECT  1.020 1.310 1.050 1.890 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 1.000 0.640 1.170 ;
        RECT  0.450 1.000 0.550 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1009 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.910 0.355 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.775 -0.330 1.200 0.330 ;
        RECT  0.665 -0.330 0.775 0.600 ;
        RECT  0.000 -0.330 0.665 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.800 2.070 1.200 2.730 ;
        RECT  0.690 1.600 0.800 2.730 ;
        RECT  0.220 2.070 0.690 2.730 ;
        RECT  0.110 1.400 0.220 2.730 ;
        RECT  0.000 2.070 0.110 2.730 ;
        END
    END VDD
END CELL91

MACRO CELL64
    CLASS CORE ;
    FOREIGN CELL64 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 0.2724 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.225 0.495 1.350 1.905 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.790 0.910 0.950 1.290 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1009 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.910 0.590 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.910 0.355 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.030 -0.330 1.400 0.330 ;
        RECT  0.920 -0.330 1.030 0.600 ;
        RECT  0.000 -0.330 0.920 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.065 2.070 1.400 2.730 ;
        RECT  0.955 1.600 1.065 2.730 ;
        RECT  0.495 2.070 0.955 2.730 ;
        RECT  0.385 1.600 0.495 2.730 ;
        RECT  0.000 2.070 0.385 2.730 ;
        END
    END VDD
END CELL64

MACRO CELL3
    CLASS CORE ;
    FOREIGN CELL3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 0.2724 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.425 0.495 1.550 1.905 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.1009 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.980 0.910 1.150 1.290 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.910 0.800 1.290 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.910 0.555 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.190 0.910 0.350 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.255 -0.330 1.600 0.330 ;
        RECT  1.145 -0.330 1.255 0.600 ;
        RECT  0.000 -0.330 1.145 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.255 2.070 1.600 2.730 ;
        RECT  1.145 1.600 1.255 2.730 ;
        RECT  0.720 2.070 1.145 2.730 ;
        RECT  0.610 1.600 0.720 2.730 ;
        RECT  0.200 2.070 0.610 2.730 ;
        RECT  0.090 1.400 0.200 2.730 ;
        RECT  0.000 2.070 0.090 2.730 ;
        END
    END VDD
END CELL3

MACRO CELL71
    CLASS CORE ;
    FOREIGN CELL71 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 0.2892 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.490 1.550 1.905 ;
        RECT  1.365 0.490 1.450 0.600 ;
        RECT  1.405 1.310 1.450 1.905 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.1009 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.995 0.910 1.150 1.290 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.910 0.795 1.290 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.1009 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.910 0.560 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.170 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.240 -0.330 1.600 0.330 ;
        RECT  1.130 -0.330 1.240 0.600 ;
        RECT  0.705 -0.330 1.130 0.330 ;
        RECT  0.595 -0.330 0.705 0.600 ;
        RECT  0.000 -0.330 0.595 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.240 2.070 1.600 2.730 ;
        RECT  1.130 1.400 1.240 2.730 ;
        RECT  0.000 2.070 1.130 2.730 ;
        END
    END VDD
END CELL71

MACRO CELL19
    CLASS CORE ;
    FOREIGN CELL19 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 0.2892 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.215 0.495 1.350 1.905 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.910 0.790 1.290 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.170 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.910 0.560 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.015 -0.330 1.400 0.330 ;
        RECT  0.905 -0.330 1.015 0.600 ;
        RECT  0.175 -0.330 0.905 0.330 ;
        RECT  0.065 -0.330 0.175 0.800 ;
        RECT  0.000 -0.330 0.065 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.015 2.070 1.400 2.730 ;
        RECT  0.905 1.400 1.015 2.730 ;
        RECT  0.000 2.070 0.905 2.730 ;
        END
    END VDD
END CELL19

MACRO CELL49
    CLASS CORE ;
    FOREIGN CELL49 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 0.1344 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.825 0.495 1.950 1.690 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.440 0.910 1.555 1.290 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.0513 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.865 0.700 0.975 0.930 ;
        RECT  0.170 0.700 0.865 0.800 ;
        RECT  0.050 0.700 0.170 1.290 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0507 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.910 1.350 1.290 ;
        RECT  1.050 1.025 1.245 1.135 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0508 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.910 0.765 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0507 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.430 0.910 0.550 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.670 -0.330 2.000 0.330 ;
        RECT  1.560 -0.330 1.670 0.600 ;
        RECT  0.000 -0.330 1.560 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.645 2.070 2.000 2.730 ;
        RECT  1.535 1.600 1.645 2.730 ;
        RECT  0.000 2.070 1.535 2.730 ;
        END
    END VDD
END CELL49

MACRO CELL42
    CLASS CORE ;
    FOREIGN CELL42 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 0.1440 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.490 1.550 1.890 ;
        RECT  1.355 0.490 1.450 0.600 ;
        RECT  1.415 1.710 1.450 1.890 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 0.890 0.285 1.000 ;
        RECT  0.050 0.890 0.150 1.290 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0506 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 1.160 1.180 1.330 ;
        RECT  1.050 0.980 1.150 1.330 ;
        RECT  0.950 0.980 1.050 1.090 ;
        RECT  0.850 0.690 0.950 1.090 ;
        RECT  0.550 0.690 0.850 0.780 ;
        RECT  0.440 0.690 0.550 0.920 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0508 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.755 1.220 0.865 1.330 ;
        RECT  0.645 0.910 0.755 1.330 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 1.110 0.555 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.180 -0.330 1.600 0.330 ;
        RECT  0.070 -0.330 0.180 0.600 ;
        RECT  0.000 -0.330 0.070 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.265 2.070 1.600 2.730 ;
        RECT  1.155 1.800 1.265 2.730 ;
        RECT  0.180 2.070 1.155 2.730 ;
        RECT  0.070 1.600 0.180 2.730 ;
        RECT  0.000 2.070 0.070 2.730 ;
        END
    END VDD
END CELL42

MACRO CELL79
    CLASS CORE ;
    FOREIGN CELL79 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 0.6720 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.150 0.510 3.260 0.890 ;
        RECT  3.150 1.310 3.260 1.890 ;
        RECT  3.050 0.710 3.150 0.890 ;
        RECT  3.050 1.310 3.150 1.490 ;
        RECT  2.750 0.710 3.050 1.490 ;
        RECT  2.640 0.510 2.750 0.890 ;
        RECT  2.640 1.310 2.750 1.890 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.2017 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.035 0.910 1.150 1.340 ;
        RECT  0.180 1.250 1.035 1.340 ;
        RECT  0.050 0.910 0.180 1.340 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2017 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.975 0.750 1.125 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.2017 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.045 0.910 2.155 1.325 ;
        RECT  1.385 1.235 2.045 1.325 ;
        RECT  1.250 0.910 1.385 1.325 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2017 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.975 1.950 1.125 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.525 -0.330 3.600 0.330 ;
        RECT  3.415 -0.330 3.525 0.800 ;
        RECT  3.005 -0.330 3.415 0.330 ;
        RECT  2.895 -0.330 3.005 0.600 ;
        RECT  2.485 -0.330 2.895 0.330 ;
        RECT  2.375 -0.330 2.485 0.600 ;
        RECT  2.270 -0.330 2.375 0.330 ;
        RECT  2.160 -0.330 2.270 0.600 ;
        RECT  1.230 -0.330 2.160 0.330 ;
        RECT  1.120 -0.330 1.230 0.600 ;
        RECT  0.190 -0.330 1.120 0.330 ;
        RECT  0.080 -0.330 0.190 0.800 ;
        RECT  0.000 -0.330 0.080 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.525 2.070 3.600 2.730 ;
        RECT  3.415 1.400 3.525 2.730 ;
        RECT  3.005 2.070 3.415 2.730 ;
        RECT  2.895 1.600 3.005 2.730 ;
        RECT  2.485 2.070 2.895 2.730 ;
        RECT  2.375 2.000 2.485 2.730 ;
        RECT  0.970 2.070 2.375 2.730 ;
        RECT  0.860 1.800 0.970 2.730 ;
        RECT  0.450 2.070 0.860 2.730 ;
        RECT  0.340 1.800 0.450 2.730 ;
        RECT  0.000 2.070 0.340 2.730 ;
        END
    END VDD
END CELL79

MACRO CELL87
    CLASS CORE ;
    FOREIGN CELL87 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 0.2856 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.490 1.550 1.905 ;
        RECT  1.365 0.490 1.450 0.600 ;
        RECT  1.405 1.310 1.450 1.905 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.960 0.910 1.150 1.200 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.170 1.290 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.910 0.555 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.910 0.790 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.240 -0.330 1.600 0.330 ;
        RECT  1.130 -0.330 1.240 0.600 ;
        RECT  0.185 -0.330 1.130 0.330 ;
        RECT  0.075 -0.330 0.185 0.600 ;
        RECT  0.000 -0.330 0.075 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.240 2.070 1.600 2.730 ;
        RECT  1.130 1.400 1.240 2.730 ;
        RECT  0.000 2.070 1.130 2.730 ;
        END
    END VDD
END CELL87

MACRO CELL85
    CLASS CORE ;
    FOREIGN CELL85 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 0.2688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.440 1.950 1.905 ;
        RECT  1.820 0.440 1.850 0.610 ;
        RECT  1.820 1.310 1.850 1.905 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.910 1.380 1.290 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.035 0.910 1.150 1.290 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.170 1.290 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.910 0.555 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.910 0.780 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.580 -0.330 2.000 0.330 ;
        RECT  1.470 -0.330 1.580 0.600 ;
        RECT  0.185 -0.330 1.470 0.330 ;
        RECT  0.075 -0.330 0.185 0.600 ;
        RECT  0.000 -0.330 0.075 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.670 2.070 2.000 2.730 ;
        RECT  1.560 2.000 1.670 2.730 ;
        RECT  1.225 2.070 1.560 2.730 ;
        RECT  1.115 1.600 1.225 2.730 ;
        RECT  0.000 2.070 1.115 2.730 ;
        END
    END VDD
END CELL85

MACRO CELL106
    CLASS CORE ;
    FOREIGN CELL106 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.2274 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.855 0.510 0.965 0.800 ;
        RECT  0.355 0.690 0.855 0.800 ;
        RECT  0.355 1.440 0.485 1.550 ;
        RECT  0.250 0.690 0.355 1.550 ;
        RECT  0.185 0.690 0.250 0.800 ;
        RECT  0.075 0.510 0.185 0.800 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.995 0.910 1.150 1.290 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.910 0.795 1.290 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.910 0.560 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.160 1.320 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.240 -0.330 1.400 0.330 ;
        RECT  1.130 -0.330 1.240 0.600 ;
        RECT  0.705 -0.330 1.130 0.330 ;
        RECT  0.595 -0.330 0.705 0.600 ;
        RECT  0.000 -0.330 0.595 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.240 2.070 1.400 2.730 ;
        RECT  1.130 1.400 1.240 2.730 ;
        RECT  0.000 2.070 1.130 2.730 ;
        END
    END VDD
END CELL106

MACRO CELL68
    CLASS CORE ;
    FOREIGN CELL68 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.4548 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.430 0.965 0.800 ;
        RECT  0.355 0.690 0.850 0.800 ;
        RECT  0.355 1.400 0.495 1.510 ;
        RECT  0.250 0.690 0.355 1.510 ;
        RECT  0.185 0.690 0.250 0.800 ;
        RECT  0.050 0.430 0.185 0.800 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.1009 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.995 0.910 1.150 1.290 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.910 0.795 1.290 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.1009 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.910 0.560 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.160 1.320 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.225 -0.330 1.400 0.330 ;
        RECT  1.115 -0.330 1.225 0.600 ;
        RECT  0.705 -0.330 1.115 0.330 ;
        RECT  0.595 -0.330 0.705 0.600 ;
        RECT  0.000 -0.330 0.595 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.225 2.070 1.400 2.730 ;
        RECT  1.115 1.400 1.225 2.730 ;
        RECT  0.000 2.070 1.115 2.730 ;
        END
    END VDD
END CELL68

MACRO CELL70
    CLASS CORE ;
    FOREIGN CELL70 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.1680 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.700 1.150 1.290 ;
        RECT  0.715 0.700 1.050 0.800 ;
        RECT  0.605 0.495 0.715 0.800 ;
        RECT  0.355 0.700 0.605 0.800 ;
        RECT  0.355 1.480 0.505 1.590 ;
        RECT  0.265 0.700 0.355 1.590 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.910 0.790 1.290 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.170 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.910 0.560 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.975 -0.330 1.200 0.330 ;
        RECT  0.865 -0.330 0.975 0.600 ;
        RECT  0.175 -0.330 0.865 0.330 ;
        RECT  0.065 -0.330 0.175 0.600 ;
        RECT  0.000 -0.330 0.065 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.975 2.070 1.200 2.730 ;
        RECT  0.865 1.400 0.975 2.730 ;
        RECT  0.000 2.070 0.865 2.730 ;
        END
    END VDD
END CELL70

MACRO CELL26
    CLASS CORE ;
    FOREIGN CELL26 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.3360 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.700 1.150 1.290 ;
        RECT  0.715 0.700 1.050 0.800 ;
        RECT  0.605 0.430 0.715 0.800 ;
        RECT  0.355 0.700 0.605 0.800 ;
        RECT  0.355 1.480 0.505 1.590 ;
        RECT  0.265 0.700 0.355 1.590 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.910 0.790 1.290 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.170 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.910 0.560 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.975 -0.330 1.200 0.330 ;
        RECT  0.865 -0.330 0.975 0.600 ;
        RECT  0.175 -0.330 0.865 0.330 ;
        RECT  0.065 -0.330 0.175 0.800 ;
        RECT  0.000 -0.330 0.065 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.975 2.070 1.200 2.730 ;
        RECT  0.865 1.400 0.975 2.730 ;
        RECT  0.000 2.070 0.865 2.730 ;
        END
    END VDD
END CELL26

MACRO CELL55
    CLASS CORE ;
    FOREIGN CELL55 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.2406 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.490 1.540 0.600 ;
        RECT  0.350 1.400 1.070 1.500 ;
        RECT  0.260 0.490 0.350 1.500 ;
        RECT  0.250 0.710 0.260 1.500 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.160 1.320 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.0514 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.440 0.710 1.550 1.290 ;
        RECT  0.765 0.710 1.440 0.800 ;
        RECT  0.650 0.710 0.765 0.940 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0508 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.910 0.555 1.290 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0511 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 1.090 0.950 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0507 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.910 1.185 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.170 -0.330 1.600 0.330 ;
        RECT  0.060 -0.330 0.170 0.600 ;
        RECT  0.000 -0.330 0.060 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.180 2.070 1.600 2.730 ;
        RECT  0.070 1.600 0.180 2.730 ;
        RECT  0.000 2.070 0.070 2.730 ;
        END
    END VDD
END CELL55

MACRO CELL13
    CLASS CORE ;
    FOREIGN CELL13 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.2418 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.560 0.490 1.890 0.600 ;
        RECT  0.355 1.400 1.450 1.510 ;
        RECT  0.450 0.490 0.560 0.800 ;
        RECT  0.355 0.710 0.450 0.800 ;
        RECT  0.250 0.710 0.355 1.510 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.0506 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.160 1.320 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.0506 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 0.910 0.560 1.290 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.0514 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.830 0.710 1.950 1.290 ;
        RECT  1.140 0.710 1.830 0.800 ;
        RECT  1.045 0.710 1.140 0.960 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0507 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 0.910 0.955 1.290 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0512 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.910 1.350 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0507 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.910 1.570 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.230 -0.330 2.000 0.330 ;
        RECT  0.120 -0.330 0.230 0.600 ;
        RECT  0.000 -0.330 0.120 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.515 2.070 2.000 2.730 ;
        RECT  0.405 1.800 0.515 2.730 ;
        RECT  0.000 2.070 0.405 2.730 ;
        END
    END VDD
END CELL13

MACRO CELL6
    CLASS CORE ;
    FOREIGN CELL6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.2274 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.690 1.350 1.510 ;
        RECT  1.220 0.690 1.250 0.800 ;
        RECT  0.810 1.400 1.250 1.510 ;
        RECT  1.110 0.510 1.220 0.800 ;
        RECT  0.180 0.690 1.110 0.800 ;
        RECT  0.070 0.510 0.180 0.800 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.910 0.555 1.290 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.170 1.290 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.910 0.770 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.910 1.155 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.700 -0.330 1.400 0.330 ;
        RECT  0.590 -0.330 0.700 0.600 ;
        RECT  0.000 -0.330 0.590 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.440 2.070 1.400 2.730 ;
        RECT  0.330 1.600 0.440 2.730 ;
        RECT  0.000 2.070 0.330 2.730 ;
        END
    END VDD
END CELL6

MACRO CELL101
    CLASS CORE ;
    FOREIGN CELL101 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.4548 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.690 1.350 1.510 ;
        RECT  1.220 0.690 1.250 0.800 ;
        RECT  0.810 1.400 1.250 1.510 ;
        RECT  1.050 0.430 1.220 0.800 ;
        RECT  0.180 0.690 1.050 0.800 ;
        RECT  0.050 0.430 0.180 0.800 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.910 0.555 1.290 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.170 1.290 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.910 0.770 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.910 1.155 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.700 -0.330 1.400 0.330 ;
        RECT  0.590 -0.330 0.700 0.600 ;
        RECT  0.000 -0.330 0.590 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.440 2.070 1.400 2.730 ;
        RECT  0.330 1.600 0.440 2.730 ;
        RECT  0.000 2.070 0.330 2.730 ;
        END
    END VDD
END CELL101

MACRO CELL21
    CLASS CORE ;
    FOREIGN CELL21 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.2448 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.855 0.495 0.965 0.800 ;
        RECT  0.350 0.700 0.855 0.800 ;
        RECT  0.350 1.400 0.745 1.510 ;
        RECT  0.250 0.700 0.350 1.510 ;
        RECT  0.185 1.400 0.250 1.510 ;
        RECT  0.050 1.400 0.185 1.800 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.960 0.910 1.150 1.200 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.880 0.160 1.290 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.910 0.555 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.910 0.790 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.225 -0.330 1.400 0.330 ;
        RECT  1.115 -0.330 1.225 0.600 ;
        RECT  0.185 -0.330 1.115 0.330 ;
        RECT  0.075 -0.330 0.185 0.600 ;
        RECT  0.000 -0.330 0.075 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.225 2.070 1.400 2.730 ;
        RECT  1.115 1.400 1.225 2.730 ;
        RECT  0.000 2.070 1.115 2.730 ;
        END
    END VDD
END CELL21

MACRO CELL4
    CLASS CORE ;
    FOREIGN CELL4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.4896 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.855 0.430 0.965 0.800 ;
        RECT  0.350 0.700 0.855 0.800 ;
        RECT  0.350 1.400 0.745 1.510 ;
        RECT  0.250 0.700 0.350 1.510 ;
        RECT  0.185 1.400 0.250 1.510 ;
        RECT  0.050 1.400 0.185 1.800 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.960 0.910 1.150 1.200 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.880 0.160 1.290 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.910 0.555 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.910 0.790 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.225 -0.330 1.400 0.330 ;
        RECT  1.115 -0.330 1.225 0.800 ;
        RECT  0.185 -0.330 1.115 0.330 ;
        RECT  0.075 -0.330 0.185 0.600 ;
        RECT  0.000 -0.330 0.075 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.225 2.070 1.400 2.730 ;
        RECT  1.115 1.400 1.225 2.730 ;
        RECT  0.000 2.070 1.115 2.730 ;
        END
    END VDD
END CELL4

MACRO CELL95
    CLASS CORE ;
    FOREIGN CELL95 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.4896 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.430 0.965 0.800 ;
        RECT  0.350 0.700 0.850 0.800 ;
        RECT  0.350 1.400 0.745 1.510 ;
        RECT  0.250 0.700 0.350 1.510 ;
        RECT  0.185 1.400 0.250 1.510 ;
        RECT  0.050 1.400 0.185 1.800 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.1009 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 0.910 1.360 1.290 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.035 0.910 1.150 1.290 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.900 0.160 1.290 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.910 0.555 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.910 0.780 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.485 -0.330 1.600 0.330 ;
        RECT  1.375 -0.330 1.485 0.600 ;
        RECT  0.185 -0.330 1.375 0.330 ;
        RECT  0.075 -0.330 0.185 0.600 ;
        RECT  0.000 -0.330 0.075 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.225 2.070 1.600 2.730 ;
        RECT  1.115 1.600 1.225 2.730 ;
        RECT  0.000 2.070 1.115 2.730 ;
        END
    END VDD
END CELL95

MACRO CELL81
    CLASS CORE ;
    FOREIGN CELL81 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.4896 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.430 0.965 0.800 ;
        RECT  0.350 0.710 0.850 0.800 ;
        RECT  0.350 1.400 0.745 1.510 ;
        RECT  0.250 0.710 0.350 1.510 ;
        RECT  0.185 1.400 0.250 1.510 ;
        RECT  0.050 1.400 0.185 1.800 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.600 0.910 1.750 1.290 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.910 1.375 1.290 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.910 1.150 1.290 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.880 0.160 1.290 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.910 0.560 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.910 0.780 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.745 -0.330 2.000 0.330 ;
        RECT  1.635 -0.330 1.745 0.600 ;
        RECT  0.185 -0.330 1.635 0.330 ;
        RECT  0.075 -0.330 0.185 0.600 ;
        RECT  0.000 -0.330 0.075 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.745 2.070 2.000 2.730 ;
        RECT  1.635 1.400 1.745 2.730 ;
        RECT  1.225 2.070 1.635 2.730 ;
        RECT  1.115 1.600 1.225 2.730 ;
        RECT  0.000 2.070 1.115 2.730 ;
        END
    END VDD
END CELL81

MACRO CELL84
    CLASS CORE ;
    FOREIGN CELL84 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 0.1344 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.625 0.510 0.750 1.800 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 1.110 0.350 1.290 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.455 -0.330 0.800 0.330 ;
        RECT  0.345 -0.330 0.455 0.600 ;
        RECT  0.000 -0.330 0.345 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.455 2.070 0.800 2.730 ;
        RECT  0.345 1.600 0.455 2.730 ;
        RECT  0.000 2.070 0.345 2.730 ;
        END
    END VDD
END CELL84

MACRO CELL73
    CLASS CORE ;
    FOREIGN CELL73 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 2.0160 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 0.510 4.170 0.890 ;
        RECT  4.050 1.310 4.170 1.890 ;
        RECT  3.650 0.710 4.050 0.890 ;
        RECT  3.650 1.310 4.050 1.490 ;
        RECT  3.540 0.510 3.650 0.890 ;
        RECT  3.540 1.310 3.650 1.890 ;
        RECT  3.150 0.710 3.540 0.890 ;
        RECT  3.150 1.310 3.540 1.490 ;
        RECT  3.050 0.510 3.150 0.890 ;
        RECT  3.050 1.310 3.150 1.890 ;
        RECT  3.025 0.510 3.050 1.890 ;
        RECT  2.610 0.710 3.025 1.490 ;
        RECT  2.550 0.510 2.610 1.890 ;
        RECT  2.500 0.510 2.550 0.890 ;
        RECT  2.500 1.310 2.550 1.890 ;
        RECT  2.090 0.710 2.500 0.890 ;
        RECT  2.090 1.310 2.500 1.490 ;
        RECT  1.980 0.510 2.090 0.890 ;
        RECT  1.980 1.310 2.090 1.890 ;
        RECT  1.565 0.710 1.980 0.890 ;
        RECT  1.565 1.310 1.980 1.490 ;
        RECT  1.450 0.510 1.565 0.890 ;
        RECT  1.450 1.310 1.565 1.890 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.4034 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 1.035 0.950 1.205 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.430 -0.330 4.600 0.330 ;
        RECT  4.320 -0.330 4.430 0.800 ;
        RECT  3.910 -0.330 4.320 0.330 ;
        RECT  3.800 -0.330 3.910 0.600 ;
        RECT  3.390 -0.330 3.800 0.330 ;
        RECT  3.280 -0.330 3.390 0.600 ;
        RECT  2.870 -0.330 3.280 0.330 ;
        RECT  2.760 -0.330 2.870 0.600 ;
        RECT  2.350 -0.330 2.760 0.330 ;
        RECT  2.240 -0.330 2.350 0.600 ;
        RECT  1.830 -0.330 2.240 0.330 ;
        RECT  1.720 -0.330 1.830 0.600 ;
        RECT  1.265 -0.330 1.720 0.330 ;
        RECT  1.155 -0.330 1.265 0.600 ;
        RECT  0.705 -0.330 1.155 0.330 ;
        RECT  0.595 -0.330 0.705 0.600 ;
        RECT  0.185 -0.330 0.595 0.330 ;
        RECT  0.075 -0.330 0.185 0.800 ;
        RECT  0.000 -0.330 0.075 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.430 2.070 4.600 2.730 ;
        RECT  4.320 1.400 4.430 2.730 ;
        RECT  3.910 2.070 4.320 2.730 ;
        RECT  3.800 1.600 3.910 2.730 ;
        RECT  3.390 2.070 3.800 2.730 ;
        RECT  3.280 1.600 3.390 2.730 ;
        RECT  2.870 2.070 3.280 2.730 ;
        RECT  2.760 1.600 2.870 2.730 ;
        RECT  2.350 2.070 2.760 2.730 ;
        RECT  2.240 1.600 2.350 2.730 ;
        RECT  1.830 2.070 2.240 2.730 ;
        RECT  1.720 1.600 1.830 2.730 ;
        RECT  1.265 2.070 1.720 2.730 ;
        RECT  1.155 1.660 1.265 2.730 ;
        RECT  0.705 2.070 1.155 2.730 ;
        RECT  0.595 1.660 0.705 2.730 ;
        RECT  0.185 2.070 0.595 2.730 ;
        RECT  0.075 1.400 0.185 2.730 ;
        RECT  0.000 2.070 0.075 2.730 ;
        END
    END VDD
END CELL73

MACRO CELL98
    CLASS CORE ;
    FOREIGN CELL98 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.800 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 2.6880 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.290 0.510 5.400 0.890 ;
        RECT  5.290 1.310 5.400 1.890 ;
        RECT  4.880 0.710 5.290 0.890 ;
        RECT  4.880 1.310 5.290 1.490 ;
        RECT  4.770 0.510 4.880 0.890 ;
        RECT  4.770 1.310 4.880 1.890 ;
        RECT  4.360 0.710 4.770 0.890 ;
        RECT  4.360 1.310 4.770 1.490 ;
        RECT  4.250 0.510 4.360 0.890 ;
        RECT  4.250 1.310 4.360 1.890 ;
        RECT  3.840 0.710 4.250 0.890 ;
        RECT  3.840 1.310 4.250 1.490 ;
        RECT  3.730 0.510 3.840 0.890 ;
        RECT  3.730 1.310 3.840 1.890 ;
        RECT  3.650 0.710 3.730 0.890 ;
        RECT  3.650 1.310 3.730 1.490 ;
        RECT  3.320 0.710 3.650 1.490 ;
        RECT  3.210 0.510 3.320 1.890 ;
        RECT  3.150 0.710 3.210 1.490 ;
        RECT  2.800 0.710 3.150 0.890 ;
        RECT  2.800 1.310 3.150 1.490 ;
        RECT  2.690 0.510 2.800 0.890 ;
        RECT  2.690 1.310 2.800 1.890 ;
        RECT  2.280 0.710 2.690 0.890 ;
        RECT  2.280 1.310 2.690 1.490 ;
        RECT  2.170 0.510 2.280 0.890 ;
        RECT  2.170 1.310 2.280 1.890 ;
        RECT  1.760 0.710 2.170 0.890 ;
        RECT  1.760 1.310 2.170 1.490 ;
        RECT  1.650 0.510 1.760 0.890 ;
        RECT  1.650 1.310 1.760 1.890 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.5042 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.035 1.150 1.205 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.660 -0.330 5.800 0.330 ;
        RECT  5.550 -0.330 5.660 0.800 ;
        RECT  5.140 -0.330 5.550 0.330 ;
        RECT  5.030 -0.330 5.140 0.600 ;
        RECT  4.620 -0.330 5.030 0.330 ;
        RECT  4.510 -0.330 4.620 0.600 ;
        RECT  4.100 -0.330 4.510 0.330 ;
        RECT  3.990 -0.330 4.100 0.600 ;
        RECT  3.580 -0.330 3.990 0.330 ;
        RECT  3.470 -0.330 3.580 0.600 ;
        RECT  3.060 -0.330 3.470 0.330 ;
        RECT  2.950 -0.330 3.060 0.600 ;
        RECT  2.540 -0.330 2.950 0.330 ;
        RECT  2.430 -0.330 2.540 0.600 ;
        RECT  2.020 -0.330 2.430 0.330 ;
        RECT  1.910 -0.330 2.020 0.600 ;
        RECT  1.500 -0.330 1.910 0.330 ;
        RECT  1.390 -0.330 1.500 0.600 ;
        RECT  0.980 -0.330 1.390 0.330 ;
        RECT  0.870 -0.330 0.980 0.600 ;
        RECT  0.460 -0.330 0.870 0.330 ;
        RECT  0.350 -0.330 0.460 0.600 ;
        RECT  0.000 -0.330 0.350 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.660 2.070 5.800 2.730 ;
        RECT  5.550 1.400 5.660 2.730 ;
        RECT  5.140 2.070 5.550 2.730 ;
        RECT  5.030 1.600 5.140 2.730 ;
        RECT  4.620 2.070 5.030 2.730 ;
        RECT  4.510 1.600 4.620 2.730 ;
        RECT  4.100 2.070 4.510 2.730 ;
        RECT  3.990 1.600 4.100 2.730 ;
        RECT  3.580 2.070 3.990 2.730 ;
        RECT  3.470 1.600 3.580 2.730 ;
        RECT  3.060 2.070 3.470 2.730 ;
        RECT  2.950 1.600 3.060 2.730 ;
        RECT  2.540 2.070 2.950 2.730 ;
        RECT  2.430 1.600 2.540 2.730 ;
        RECT  2.020 2.070 2.430 2.730 ;
        RECT  1.910 1.600 2.020 2.730 ;
        RECT  1.500 2.070 1.910 2.730 ;
        RECT  1.390 1.690 1.500 2.730 ;
        RECT  0.980 2.070 1.390 2.730 ;
        RECT  0.870 1.690 0.980 2.730 ;
        RECT  0.460 2.070 0.870 2.730 ;
        RECT  0.350 1.690 0.460 2.730 ;
        RECT  0.000 2.070 0.350 2.730 ;
        END
    END VDD
END CELL98

MACRO CELL38
    CLASS CORE ;
    FOREIGN CELL38 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 0.2688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.625 0.510 0.750 1.890 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0582 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 1.110 0.350 1.290 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.455 -0.330 0.800 0.330 ;
        RECT  0.345 -0.330 0.455 0.600 ;
        RECT  0.000 -0.330 0.345 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.455 2.070 0.800 2.730 ;
        RECT  0.345 1.600 0.455 2.730 ;
        RECT  0.000 2.070 0.345 2.730 ;
        END
    END VDD
END CELL38

MACRO CELL67
    CLASS CORE ;
    FOREIGN CELL67 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 0.3360 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.510 0.775 1.890 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.350 1.125 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.030 -0.330 1.200 0.330 ;
        RECT  0.920 -0.330 1.030 0.800 ;
        RECT  0.485 -0.330 0.920 0.330 ;
        RECT  0.375 -0.330 0.485 0.600 ;
        RECT  0.000 -0.330 0.375 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.030 2.070 1.200 2.730 ;
        RECT  0.920 1.400 1.030 2.730 ;
        RECT  0.485 2.070 0.920 2.730 ;
        RECT  0.375 1.600 0.485 2.730 ;
        RECT  0.000 2.070 0.375 2.730 ;
        END
    END VDD
END CELL67

MACRO CELL48
    CLASS CORE ;
    FOREIGN CELL48 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 0.6720 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.510 1.570 0.890 ;
        RECT  1.450 1.310 1.570 1.890 ;
        RECT  1.150 0.710 1.450 1.490 ;
        RECT  1.050 0.710 1.150 0.890 ;
        RECT  1.050 1.310 1.150 1.490 ;
        RECT  0.940 0.510 1.050 0.890 ;
        RECT  0.940 1.310 1.050 1.890 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.2017 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.910 0.550 1.290 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.835 -0.330 2.000 0.330 ;
        RECT  1.725 -0.330 1.835 0.800 ;
        RECT  1.315 -0.330 1.725 0.330 ;
        RECT  1.205 -0.330 1.315 0.600 ;
        RECT  0.760 -0.330 1.205 0.330 ;
        RECT  0.650 -0.330 0.760 0.600 ;
        RECT  0.240 -0.330 0.650 0.330 ;
        RECT  0.130 -0.330 0.240 0.800 ;
        RECT  0.000 -0.330 0.130 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.835 2.070 2.000 2.730 ;
        RECT  1.725 1.400 1.835 2.730 ;
        RECT  1.315 2.070 1.725 2.730 ;
        RECT  1.205 1.600 1.315 2.730 ;
        RECT  0.760 2.070 1.205 2.730 ;
        RECT  0.650 1.600 0.760 2.730 ;
        RECT  0.240 2.070 0.650 2.730 ;
        RECT  0.130 1.400 0.240 2.730 ;
        RECT  0.000 2.070 0.130 2.730 ;
        END
    END VDD
END CELL48

MACRO CELL45
    CLASS CORE ;
    FOREIGN CELL45 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 1.0080 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.925 0.510 2.035 0.890 ;
        RECT  1.925 1.310 2.035 1.890 ;
        RECT  1.650 0.710 1.925 0.890 ;
        RECT  1.650 1.310 1.925 1.490 ;
        RECT  1.515 0.710 1.650 1.490 ;
        RECT  1.405 0.510 1.515 1.890 ;
        RECT  1.350 0.710 1.405 1.490 ;
        RECT  0.995 0.710 1.350 0.890 ;
        RECT  0.995 1.310 1.350 1.490 ;
        RECT  0.885 0.510 0.995 0.890 ;
        RECT  0.885 1.310 0.995 1.890 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.2017 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.910 0.550 1.290 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.295 -0.330 2.400 0.330 ;
        RECT  2.185 -0.330 2.295 0.800 ;
        RECT  1.775 -0.330 2.185 0.330 ;
        RECT  1.665 -0.330 1.775 0.600 ;
        RECT  1.255 -0.330 1.665 0.330 ;
        RECT  1.145 -0.330 1.255 0.600 ;
        RECT  0.735 -0.330 1.145 0.330 ;
        RECT  0.625 -0.330 0.735 0.600 ;
        RECT  0.215 -0.330 0.625 0.330 ;
        RECT  0.105 -0.330 0.215 0.800 ;
        RECT  0.000 -0.330 0.105 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.295 2.070 2.400 2.730 ;
        RECT  2.185 1.400 2.295 2.730 ;
        RECT  1.775 2.070 2.185 2.730 ;
        RECT  1.665 1.600 1.775 2.730 ;
        RECT  1.255 2.070 1.665 2.730 ;
        RECT  1.145 1.600 1.255 2.730 ;
        RECT  0.735 2.070 1.145 2.730 ;
        RECT  0.625 1.600 0.735 2.730 ;
        RECT  0.215 2.070 0.625 2.730 ;
        RECT  0.105 1.400 0.215 2.730 ;
        RECT  0.000 2.070 0.105 2.730 ;
        END
    END VDD
END CELL45

MACRO CELL16
    CLASS CORE ;
    FOREIGN CELL16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 1.3440 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.700 0.510 2.810 0.890 ;
        RECT  2.700 1.310 2.810 1.890 ;
        RECT  2.290 0.710 2.700 0.890 ;
        RECT  2.290 1.310 2.700 1.490 ;
        RECT  2.250 0.510 2.290 0.890 ;
        RECT  2.250 1.310 2.290 1.890 ;
        RECT  2.180 0.510 2.250 1.890 ;
        RECT  1.765 0.710 2.180 1.490 ;
        RECT  1.750 0.510 1.765 1.890 ;
        RECT  1.650 0.510 1.750 0.890 ;
        RECT  1.650 1.310 1.750 1.890 ;
        RECT  1.250 0.710 1.650 0.890 ;
        RECT  1.250 1.310 1.650 1.490 ;
        RECT  1.140 0.510 1.250 0.890 ;
        RECT  1.140 1.310 1.250 1.890 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.3026 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 1.030 0.750 1.270 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.070 -0.330 3.200 0.330 ;
        RECT  2.960 -0.330 3.070 0.800 ;
        RECT  2.550 -0.330 2.960 0.330 ;
        RECT  2.440 -0.330 2.550 0.600 ;
        RECT  2.030 -0.330 2.440 0.330 ;
        RECT  1.920 -0.330 2.030 0.600 ;
        RECT  1.510 -0.330 1.920 0.330 ;
        RECT  1.400 -0.330 1.510 0.600 ;
        RECT  0.990 -0.330 1.400 0.330 ;
        RECT  0.880 -0.330 0.990 0.600 ;
        RECT  0.470 -0.330 0.880 0.330 ;
        RECT  0.360 -0.330 0.470 0.600 ;
        RECT  0.000 -0.330 0.360 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.070 2.070 3.200 2.730 ;
        RECT  2.960 1.400 3.070 2.730 ;
        RECT  2.550 2.070 2.960 2.730 ;
        RECT  2.440 1.600 2.550 2.730 ;
        RECT  2.030 2.070 2.440 2.730 ;
        RECT  1.920 1.600 2.030 2.730 ;
        RECT  1.510 2.070 1.920 2.730 ;
        RECT  1.400 1.600 1.510 2.730 ;
        RECT  0.990 2.070 1.400 2.730 ;
        RECT  0.880 1.610 0.990 2.730 ;
        RECT  0.470 2.070 0.880 2.730 ;
        RECT  0.360 1.610 0.470 2.730 ;
        RECT  0.000 2.070 0.360 2.730 ;
        END
    END VDD
END CELL16

MACRO CELL2
    CLASS CORE ;
    FOREIGN CELL2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 0.1314 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.455 1.150 1.800 ;
        RECT  0.980 0.455 1.050 0.635 ;
        RECT  0.980 1.400 1.050 1.800 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 1.000 0.640 1.230 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.910 0.355 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.775 -0.330 1.200 0.330 ;
        RECT  0.665 -0.330 0.775 0.575 ;
        RECT  0.000 -0.330 0.665 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.800 2.070 1.200 2.730 ;
        RECT  0.690 1.600 0.800 2.730 ;
        RECT  0.220 2.070 0.690 2.730 ;
        RECT  0.110 1.400 0.220 2.730 ;
        RECT  0.000 2.070 0.110 2.730 ;
        END
    END VDD
END CELL2

MACRO CELL82
    CLASS CORE ;
    FOREIGN CELL82 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 0.2484 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.465 1.150 1.890 ;
        RECT  0.980 0.465 1.050 0.845 ;
        RECT  1.020 1.310 1.050 1.890 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0512 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 1.000 0.640 1.230 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.910 0.355 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.775 -0.330 1.200 0.330 ;
        RECT  0.665 -0.330 0.775 0.600 ;
        RECT  0.000 -0.330 0.665 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.820 2.070 1.200 2.730 ;
        RECT  0.710 1.800 0.820 2.730 ;
        RECT  0.225 2.070 0.710 2.730 ;
        RECT  0.105 1.600 0.225 2.730 ;
        RECT  0.000 2.070 0.105 2.730 ;
        END
    END VDD
END CELL82

MACRO CELL77
    CLASS CORE ;
    FOREIGN CELL77 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 2.3070 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.510 4.860 0.690 ;
        RECT  4.750 1.110 4.860 1.890 ;
        RECT  4.350 1.110 4.750 1.290 ;
        RECT  4.230 1.110 4.350 1.890 ;
        RECT  3.820 1.110 4.230 1.290 ;
        RECT  3.710 1.110 3.820 1.890 ;
        RECT  3.450 1.110 3.710 1.290 ;
        RECT  3.300 0.510 3.450 1.290 ;
        RECT  3.190 0.510 3.300 1.890 ;
        RECT  2.950 0.510 3.190 1.290 ;
        RECT  1.630 0.510 2.950 0.690 ;
        RECT  2.780 1.110 2.950 1.290 ;
        RECT  2.670 1.110 2.780 1.890 ;
        RECT  2.260 1.110 2.670 1.290 ;
        RECT  2.150 1.110 2.260 1.890 ;
        RECT  1.750 1.110 2.150 1.290 ;
        RECT  1.630 1.110 1.750 1.890 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.4178 ;
        ANTENNADIFFAREA 0.0660 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.190 1.030 1.150 1.210 ;
        RECT  0.050 0.510 0.190 1.210 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.120 -0.330 5.200 0.330 ;
        RECT  5.010 -0.330 5.120 0.600 ;
        RECT  1.480 -0.330 5.010 0.330 ;
        RECT  1.370 -0.330 1.480 0.600 ;
        RECT  1.255 -0.330 1.370 0.330 ;
        RECT  1.145 -0.330 1.255 0.600 ;
        RECT  0.735 -0.330 1.145 0.330 ;
        RECT  0.625 -0.330 0.735 0.600 ;
        RECT  0.000 -0.330 0.625 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.120 2.070 5.200 2.730 ;
        RECT  5.010 1.400 5.120 2.730 ;
        RECT  4.600 2.070 5.010 2.730 ;
        RECT  4.490 1.400 4.600 2.730 ;
        RECT  4.080 2.070 4.490 2.730 ;
        RECT  3.970 1.400 4.080 2.730 ;
        RECT  3.560 2.070 3.970 2.730 ;
        RECT  3.430 1.400 3.560 2.730 ;
        RECT  3.040 2.070 3.430 2.730 ;
        RECT  2.930 1.400 3.040 2.730 ;
        RECT  2.520 2.070 2.930 2.730 ;
        RECT  2.410 1.400 2.520 2.730 ;
        RECT  2.000 2.070 2.410 2.730 ;
        RECT  1.890 1.400 2.000 2.730 ;
        RECT  1.480 2.070 1.890 2.730 ;
        RECT  1.370 1.695 1.480 2.730 ;
        RECT  0.960 2.070 1.370 2.730 ;
        RECT  0.850 1.695 0.960 2.730 ;
        RECT  0.440 2.070 0.850 2.730 ;
        RECT  0.330 1.695 0.440 2.730 ;
        RECT  0.000 2.070 0.330 2.730 ;
        END
    END VDD
END CELL77

MACRO CELL69
    CLASS CORE ;
    FOREIGN CELL69 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 0.2336 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.625 0.510 0.750 1.890 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.0876 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.350 1.090 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.455 -0.330 0.800 0.330 ;
        RECT  0.345 -0.330 0.455 0.600 ;
        RECT  0.000 -0.330 0.345 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.455 2.070 0.800 2.730 ;
        RECT  0.345 1.600 0.455 2.730 ;
        RECT  0.000 2.070 0.345 2.730 ;
        END
    END VDD
END CELL69

MACRO CELL61
    CLASS CORE ;
    FOREIGN CELL61 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 2.9460 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.450 0.510 6.350 0.690 ;
        RECT  6.200 1.110 6.350 1.890 ;
        RECT  5.790 1.110 6.200 1.290 ;
        RECT  5.680 1.110 5.790 1.890 ;
        RECT  5.270 1.110 5.680 1.290 ;
        RECT  5.160 1.110 5.270 1.890 ;
        RECT  4.750 1.110 5.160 1.290 ;
        RECT  4.640 1.110 4.750 1.890 ;
        RECT  4.450 1.110 4.640 1.290 ;
        RECT  4.230 0.510 4.450 1.290 ;
        RECT  4.120 0.510 4.230 1.890 ;
        RECT  3.950 0.510 4.120 1.290 ;
        RECT  2.040 0.510 3.950 0.690 ;
        RECT  3.710 1.110 3.950 1.290 ;
        RECT  3.600 1.110 3.710 1.890 ;
        RECT  3.190 1.110 3.600 1.290 ;
        RECT  3.080 1.110 3.190 1.890 ;
        RECT  2.670 1.110 3.080 1.290 ;
        RECT  2.560 1.110 2.670 1.890 ;
        RECT  2.150 1.110 2.560 1.290 ;
        RECT  2.040 1.110 2.150 1.890 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.5186 ;
        ANTENNADIFFAREA 0.0660 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.190 1.030 1.550 1.210 ;
        RECT  0.050 0.510 0.190 1.210 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.890 -0.330 6.400 0.330 ;
        RECT  1.780 -0.330 1.890 0.600 ;
        RECT  1.500 -0.330 1.780 0.330 ;
        RECT  1.390 -0.330 1.500 0.600 ;
        RECT  0.980 -0.330 1.390 0.330 ;
        RECT  0.870 -0.330 0.980 0.600 ;
        RECT  0.460 -0.330 0.870 0.330 ;
        RECT  0.350 -0.330 0.460 0.800 ;
        RECT  0.000 -0.330 0.350 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.050 2.070 6.400 2.730 ;
        RECT  5.940 1.400 6.050 2.730 ;
        RECT  5.530 2.070 5.940 2.730 ;
        RECT  5.420 1.400 5.530 2.730 ;
        RECT  5.010 2.070 5.420 2.730 ;
        RECT  4.900 1.400 5.010 2.730 ;
        RECT  4.490 2.070 4.900 2.730 ;
        RECT  4.380 1.400 4.490 2.730 ;
        RECT  3.970 2.070 4.380 2.730 ;
        RECT  3.860 1.400 3.970 2.730 ;
        RECT  3.450 2.070 3.860 2.730 ;
        RECT  3.340 1.400 3.450 2.730 ;
        RECT  2.930 2.070 3.340 2.730 ;
        RECT  2.820 1.400 2.930 2.730 ;
        RECT  2.410 2.070 2.820 2.730 ;
        RECT  2.300 1.400 2.410 2.730 ;
        RECT  1.860 2.070 2.300 2.730 ;
        RECT  1.750 1.800 1.860 2.730 ;
        RECT  1.310 2.070 1.750 2.730 ;
        RECT  1.200 1.800 1.310 2.730 ;
        RECT  0.790 2.070 1.200 2.730 ;
        RECT  0.680 1.800 0.790 2.730 ;
        RECT  0.270 2.070 0.680 2.730 ;
        RECT  0.160 1.400 0.270 2.730 ;
        RECT  0.000 2.070 0.160 2.730 ;
        END
    END VDD
END CELL61

MACRO CELL89
    CLASS CORE ;
    FOREIGN CELL89 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 3.3460 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.850 0.510 7.150 0.690 ;
        RECT  7.005 1.110 7.150 1.890 ;
        RECT  6.595 1.110 7.005 1.290 ;
        RECT  6.485 1.110 6.595 1.890 ;
        RECT  6.075 1.110 6.485 1.290 ;
        RECT  5.965 1.110 6.075 1.890 ;
        RECT  5.555 1.110 5.965 1.290 ;
        RECT  5.445 1.110 5.555 1.890 ;
        RECT  5.035 1.110 5.445 1.290 ;
        RECT  4.925 1.110 5.035 1.890 ;
        RECT  4.850 1.110 4.925 1.290 ;
        RECT  4.550 0.510 4.850 1.290 ;
        RECT  4.405 0.510 4.550 1.890 ;
        RECT  4.350 0.510 4.405 1.290 ;
        RECT  2.325 0.510 4.350 0.690 ;
        RECT  3.995 1.110 4.350 1.290 ;
        RECT  3.885 1.110 3.995 1.890 ;
        RECT  3.475 1.110 3.885 1.290 ;
        RECT  3.365 1.110 3.475 1.890 ;
        RECT  2.955 1.110 3.365 1.290 ;
        RECT  2.845 1.110 2.955 1.890 ;
        RECT  2.435 1.110 2.845 1.290 ;
        RECT  2.325 1.110 2.435 1.890 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.6133 ;
        ANTENNADIFFAREA 0.0660 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.190 1.030 1.645 1.210 ;
        RECT  0.050 0.510 0.190 1.210 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.375 -0.330 7.600 0.330 ;
        RECT  7.265 -0.330 7.375 0.600 ;
        RECT  2.175 -0.330 7.265 0.330 ;
        RECT  2.065 -0.330 2.175 0.570 ;
        RECT  1.765 -0.330 2.065 0.330 ;
        RECT  1.655 -0.330 1.765 0.570 ;
        RECT  1.245 -0.330 1.655 0.330 ;
        RECT  1.135 -0.330 1.245 0.570 ;
        RECT  0.725 -0.330 1.135 0.330 ;
        RECT  0.615 -0.330 0.725 0.570 ;
        RECT  0.000 -0.330 0.615 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.375 2.070 7.600 2.730 ;
        RECT  7.265 1.400 7.375 2.730 ;
        RECT  6.855 2.070 7.265 2.730 ;
        RECT  6.745 1.400 6.855 2.730 ;
        RECT  6.335 2.070 6.745 2.730 ;
        RECT  6.225 1.400 6.335 2.730 ;
        RECT  5.815 2.070 6.225 2.730 ;
        RECT  5.705 1.400 5.815 2.730 ;
        RECT  5.295 2.070 5.705 2.730 ;
        RECT  5.185 1.400 5.295 2.730 ;
        RECT  4.775 2.070 5.185 2.730 ;
        RECT  4.665 1.400 4.775 2.730 ;
        RECT  4.255 2.070 4.665 2.730 ;
        RECT  4.145 1.400 4.255 2.730 ;
        RECT  3.735 2.070 4.145 2.730 ;
        RECT  3.625 1.400 3.735 2.730 ;
        RECT  3.215 2.070 3.625 2.730 ;
        RECT  3.105 1.400 3.215 2.730 ;
        RECT  2.695 2.070 3.105 2.730 ;
        RECT  2.585 1.400 2.695 2.730 ;
        RECT  2.105 2.070 2.585 2.730 ;
        RECT  1.995 1.800 2.105 2.730 ;
        RECT  1.515 2.070 1.995 2.730 ;
        RECT  1.405 1.800 1.515 2.730 ;
        RECT  0.995 2.070 1.405 2.730 ;
        RECT  0.885 1.800 0.995 2.730 ;
        RECT  0.475 2.070 0.885 2.730 ;
        RECT  0.365 1.800 0.475 2.730 ;
        RECT  0.000 2.070 0.365 2.730 ;
        END
    END VDD
END CELL89

MACRO CELL39
    CLASS CORE ;
    FOREIGN CELL39 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 1.1680 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.510 2.810 0.690 ;
        RECT  2.700 1.310 2.810 1.890 ;
        RECT  2.290 1.310 2.700 1.490 ;
        RECT  2.250 1.310 2.290 1.890 ;
        RECT  2.180 0.510 2.250 1.890 ;
        RECT  1.770 0.510 2.180 1.490 ;
        RECT  1.750 0.510 1.770 1.890 ;
        RECT  1.140 0.510 1.750 0.690 ;
        RECT  1.650 1.310 1.750 1.890 ;
        RECT  1.250 1.310 1.650 1.490 ;
        RECT  1.140 1.310 1.250 1.890 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.2593 ;
        ANTENNADIFFAREA 0.0660 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.190 1.030 0.750 1.210 ;
        RECT  0.050 0.510 0.190 1.210 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.070 -0.330 3.200 0.330 ;
        RECT  2.960 -0.330 3.070 0.600 ;
        RECT  0.990 -0.330 2.960 0.330 ;
        RECT  0.880 -0.330 0.990 0.600 ;
        RECT  0.470 -0.330 0.880 0.330 ;
        RECT  0.360 -0.330 0.470 0.800 ;
        RECT  0.000 -0.330 0.360 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.070 2.070 3.200 2.730 ;
        RECT  2.960 1.400 3.070 2.730 ;
        RECT  2.550 2.070 2.960 2.730 ;
        RECT  2.430 1.600 2.550 2.730 ;
        RECT  2.030 2.070 2.430 2.730 ;
        RECT  1.920 1.600 2.030 2.730 ;
        RECT  1.510 2.070 1.920 2.730 ;
        RECT  1.400 1.600 1.510 2.730 ;
        RECT  0.990 2.070 1.400 2.730 ;
        RECT  0.880 1.610 0.990 2.730 ;
        RECT  0.470 2.070 0.880 2.730 ;
        RECT  0.360 1.610 0.470 2.730 ;
        RECT  0.000 2.070 0.360 2.730 ;
        END
    END VDD
END CELL39

MACRO CELL78
    CLASS CORE ;
    FOREIGN CELL78 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 2.400 ;
    SYMMETRY x y ;
    PIN TE
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.170 1.290 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.5840 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 0.510 4.065 0.890 ;
        RECT  4.050 1.310 4.065 1.890 ;
        RECT  3.955 0.510 4.050 1.890 ;
        RECT  3.750 0.710 3.955 1.490 ;
        RECT  3.550 0.710 3.750 0.890 ;
        RECT  3.550 1.310 3.750 1.490 ;
        RECT  3.435 0.510 3.550 0.890 ;
        RECT  3.435 1.310 3.550 1.890 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.910 0.555 1.290 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.1265 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 1.110 2.750 1.290 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.325 -0.330 4.400 0.330 ;
        RECT  4.215 -0.330 4.325 0.800 ;
        RECT  3.805 -0.330 4.215 0.330 ;
        RECT  3.695 -0.330 3.805 0.600 ;
        RECT  3.285 -0.330 3.695 0.330 ;
        RECT  3.175 -0.330 3.285 0.800 ;
        RECT  1.565 -0.330 3.175 0.330 ;
        RECT  1.455 -0.330 1.565 0.600 ;
        RECT  0.445 -0.330 1.455 0.330 ;
        RECT  0.335 -0.330 0.445 0.600 ;
        RECT  0.000 -0.330 0.335 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.325 2.070 4.400 2.730 ;
        RECT  4.215 1.400 4.325 2.730 ;
        RECT  3.805 2.070 4.215 2.730 ;
        RECT  3.695 1.600 3.805 2.730 ;
        RECT  3.285 2.070 3.695 2.730 ;
        RECT  3.175 1.400 3.285 2.730 ;
        RECT  2.275 2.070 3.175 2.730 ;
        RECT  2.165 1.600 2.275 2.730 ;
        RECT  1.530 2.070 2.165 2.730 ;
        RECT  1.420 1.800 1.530 2.730 ;
        RECT  0.185 2.070 1.420 2.730 ;
        RECT  0.075 1.400 0.185 2.730 ;
        RECT  0.000 2.070 0.075 2.730 ;
        END
    END VDD
END CELL78

MACRO CELL83
    CLASS CORE ;
    FOREIGN CELL83 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.600 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.1484 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.600 0.550 1.800 ;
        RECT  0.375 0.600 0.450 0.800 ;
        RECT  0.375 1.400 0.450 1.800 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.0438 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 1.000 0.350 1.210 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.225 -0.330 0.600 0.330 ;
        RECT  0.115 -0.330 0.225 0.800 ;
        RECT  0.000 -0.330 0.115 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.225 2.070 0.600 2.730 ;
        RECT  0.115 1.400 0.225 2.730 ;
        RECT  0.000 2.070 0.115 2.730 ;
        END
    END VDD
END CELL83

MACRO CELL76
    CLASS CORE ;
    FOREIGN CELL76 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.2920 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.710 0.550 1.490 ;
        RECT  0.450 0.510 0.455 1.890 ;
        RECT  0.345 0.510 0.450 0.890 ;
        RECT  0.345 1.310 0.450 1.890 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.1752 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.160 1.000 0.245 1.170 ;
        RECT  0.050 1.000 0.160 1.290 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.715 -0.330 0.800 0.330 ;
        RECT  0.605 -0.330 0.715 0.600 ;
        RECT  0.195 -0.330 0.605 0.330 ;
        RECT  0.085 -0.330 0.195 0.600 ;
        RECT  0.000 -0.330 0.085 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.715 2.070 0.800 2.730 ;
        RECT  0.605 1.600 0.715 2.730 ;
        RECT  0.195 2.070 0.605 2.730 ;
        RECT  0.085 1.400 0.195 2.730 ;
        RECT  0.000 2.070 0.085 2.730 ;
        END
    END VDD
END CELL76

MACRO CELL23
    CLASS CORE ;
    FOREIGN CELL23 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.0905 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.600 0.750 1.490 ;
        RECT  0.605 0.600 0.650 0.800 ;
        RECT  0.455 1.400 0.650 1.490 ;
        RECT  0.345 1.400 0.455 1.970 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0294 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.180 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0294 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.910 0.550 1.300 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.195 -0.330 0.800 0.330 ;
        RECT  0.085 -0.330 0.195 0.800 ;
        RECT  0.000 -0.330 0.085 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.715 2.070 0.800 2.730 ;
        RECT  0.605 1.800 0.715 2.730 ;
        RECT  0.195 2.070 0.605 2.730 ;
        RECT  0.085 1.800 0.195 2.730 ;
        RECT  0.000 2.070 0.085 2.730 ;
        END
    END VDD
END CELL23

MACRO CELL51
    CLASS CORE ;
    FOREIGN CELL51 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 0.2688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.510 2.350 1.890 ;
        RECT  2.220 0.510 2.250 0.890 ;
        RECT  2.220 1.310 2.250 1.890 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.230 0.910 0.350 1.290 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.070 -0.330 2.400 0.330 ;
        RECT  1.960 -0.330 2.070 0.830 ;
        RECT  0.440 -0.330 1.960 0.330 ;
        RECT  0.330 -0.330 0.440 0.610 ;
        RECT  0.000 -0.330 0.330 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.070 2.070 2.400 2.730 ;
        RECT  1.960 1.400 2.070 2.730 ;
        RECT  0.440 2.070 1.960 2.730 ;
        RECT  0.330 1.650 0.440 2.730 ;
        RECT  0.000 2.070 0.330 2.730 ;
        END
    END VDD
END CELL51

MACRO CELL34
    CLASS CORE ;
    FOREIGN CELL34 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY x y ;
    PIN QN
        ANTENNADIFFAREA 0.3360 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.465 0.710 4.550 1.490 ;
        RECT  4.450 0.510 4.465 1.890 ;
        RECT  4.355 0.510 4.450 0.890 ;
        RECT  4.355 1.310 4.450 1.890 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3360 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.835 0.710 3.950 1.890 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0960 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 1.025 1.365 1.135 ;
        RECT  1.050 1.025 1.150 1.490 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0517 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.045 0.910 0.185 1.290 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.725 -0.330 4.800 0.330 ;
        RECT  4.615 -0.330 4.725 0.600 ;
        RECT  0.935 -0.330 4.615 0.330 ;
        RECT  0.825 -0.330 0.935 0.600 ;
        RECT  0.000 -0.330 0.825 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.725 2.070 4.800 2.730 ;
        RECT  4.615 1.600 4.725 2.730 ;
        RECT  4.205 2.070 4.615 2.730 ;
        RECT  4.095 1.400 4.205 2.730 ;
        RECT  3.665 2.070 4.095 2.730 ;
        RECT  3.555 1.800 3.665 2.730 ;
        RECT  3.125 2.070 3.555 2.730 ;
        RECT  3.015 1.800 3.125 2.730 ;
        RECT  0.000 2.070 3.015 2.730 ;
        END
    END VDD
END CELL34

MACRO CELL28
    CLASS CORE ;
    FOREIGN CELL28 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 2.400 ;
    SYMMETRY x y ;
    PIN QN
        ANTENNADIFFAREA 0.3360 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.850 0.745 3.950 1.545 ;
        RECT  3.615 0.745 3.850 0.855 ;
        RECT  3.615 1.435 3.850 1.545 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3360 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.865 0.710 4.950 1.490 ;
        RECT  4.850 0.510 4.865 1.890 ;
        RECT  4.755 0.510 4.850 0.890 ;
        RECT  4.755 1.310 4.850 1.890 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.900 1.360 1.290 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0517 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.180 1.290 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.845 0.900 0.955 1.290 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.125 -0.330 5.200 0.330 ;
        RECT  5.015 -0.330 5.125 0.600 ;
        RECT  4.605 -0.330 5.015 0.330 ;
        RECT  4.495 -0.330 4.605 0.600 ;
        RECT  0.000 -0.330 4.495 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.125 2.070 5.200 2.730 ;
        RECT  5.015 1.600 5.125 2.730 ;
        RECT  4.605 2.070 5.015 2.730 ;
        RECT  4.495 1.600 4.605 2.730 ;
        RECT  4.090 2.070 4.495 2.730 ;
        RECT  3.920 1.850 4.090 2.730 ;
        RECT  3.545 2.070 3.920 2.730 ;
        RECT  3.375 1.850 3.545 2.730 ;
        RECT  2.360 2.070 3.375 2.730 ;
        RECT  2.250 1.600 2.360 2.730 ;
        RECT  1.220 2.070 2.250 2.730 ;
        RECT  1.110 1.800 1.220 2.730 ;
        RECT  0.000 2.070 1.110 2.730 ;
        END
    END VDD
END CELL28

MACRO CELL31
    CLASS CORE ;
    FOREIGN CELL31 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 2.400 ;
    SYMMETRY x y ;
    PIN Q
        ANTENNADIFFAREA 0.2688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.050 0.510 4.150 1.890 ;
        RECT  4.015 0.510 4.050 0.890 ;
        RECT  4.015 1.310 4.050 1.890 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0900 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.910 1.350 1.290 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0517 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.170 1.290 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.0900 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.910 1.030 1.165 ;
        RECT  0.850 0.910 0.950 1.290 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.865 -0.330 4.200 0.330 ;
        RECT  3.755 -0.330 3.865 0.600 ;
        RECT  3.280 -0.330 3.755 0.330 ;
        RECT  3.170 -0.330 3.280 0.690 ;
        RECT  0.935 -0.330 3.170 0.330 ;
        RECT  0.825 -0.330 0.935 0.600 ;
        RECT  0.000 -0.330 0.825 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.865 2.070 4.200 2.730 ;
        RECT  3.755 1.800 3.865 2.730 ;
        RECT  3.345 2.070 3.755 2.730 ;
        RECT  3.235 1.580 3.345 2.730 ;
        RECT  2.315 2.070 3.235 2.730 ;
        RECT  2.205 1.600 2.315 2.730 ;
        RECT  1.250 2.070 2.205 2.730 ;
        RECT  1.080 1.850 1.250 2.730 ;
        RECT  0.000 2.070 1.080 2.730 ;
        END
    END VDD
END CELL31

MACRO CELL60
    CLASS CORE ;
    FOREIGN CELL60 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 2.400 ;
    SYMMETRY x y ;
    PIN SN
        ANTENNAGATEAREA 0.0512 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.910 1.020 1.165 ;
        RECT  0.850 0.910 0.950 1.290 ;
        END
    END SN
    PIN QN
        ANTENNADIFFAREA 0.3360 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.250 0.710 5.350 1.490 ;
        RECT  5.220 0.710 5.250 0.890 ;
        RECT  5.220 1.310 5.250 1.490 ;
        RECT  5.110 0.510 5.220 0.890 ;
        RECT  5.110 1.310 5.220 1.890 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3360 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.700 0.710 4.750 1.490 ;
        RECT  4.650 0.710 4.700 1.890 ;
        RECT  4.590 0.710 4.650 0.890 ;
        RECT  4.590 1.310 4.650 1.890 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.1009 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.430 0.910 1.550 1.290 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0517 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 1.000 0.280 1.170 ;
        RECT  0.050 0.910 0.150 1.290 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.480 -0.330 5.600 0.330 ;
        RECT  5.370 -0.330 5.480 0.600 ;
        RECT  0.000 -0.330 5.370 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.480 2.070 5.600 2.730 ;
        RECT  5.370 1.600 5.480 2.730 ;
        RECT  4.965 2.070 5.370 2.730 ;
        RECT  4.835 1.600 4.965 2.730 ;
        RECT  4.440 2.070 4.835 2.730 ;
        RECT  4.330 1.400 4.440 2.730 ;
        RECT  3.920 2.070 4.330 2.730 ;
        RECT  3.810 1.800 3.920 2.730 ;
        RECT  2.820 2.070 3.810 2.730 ;
        RECT  2.650 1.455 2.820 2.730 ;
        RECT  0.000 2.070 2.650 2.730 ;
        END
    END VDD
END CELL60

MACRO CELL17
    CLASS CORE ;
    FOREIGN CELL17 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 2.400 ;
    SYMMETRY x y ;
    PIN Q
        ANTENNADIFFAREA 0.2688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.625 0.495 3.750 1.905 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.0960 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 1.025 1.375 1.135 ;
        RECT  1.050 1.025 1.150 1.490 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0517 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.180 1.290 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.990 -0.330 3.800 0.330 ;
        RECT  2.880 -0.330 2.990 0.600 ;
        RECT  0.935 -0.330 2.880 0.330 ;
        RECT  0.825 -0.330 0.935 0.600 ;
        RECT  0.000 -0.330 0.825 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.070 3.800 2.730 ;
        END
    END VDD
END CELL17

MACRO CELL104
    CLASS CORE ;
    FOREIGN CELL104 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 2.400 ;
    SYMMETRY x y ;
    PIN QN
        ANTENNADIFFAREA 0.2772 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.420 0.495 5.550 1.905 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.2940 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.050 0.710 5.150 1.490 ;
        RECT  4.840 0.710 5.050 0.890 ;
        RECT  4.840 1.310 5.050 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.1334 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.910 0.360 1.300 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0772 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.995 0.590 1.165 ;
        RECT  0.450 0.710 0.550 1.165 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0511 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 0.910 1.750 1.165 ;
        RECT  1.450 0.910 1.640 1.090 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.210 -0.330 5.600 0.330 ;
        RECT  3.100 -0.330 3.210 0.810 ;
        RECT  0.485 -0.330 3.100 0.330 ;
        RECT  0.315 -0.330 0.485 0.600 ;
        RECT  0.000 -0.330 0.315 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.230 2.070 5.600 2.730 ;
        RECT  3.060 1.800 3.230 2.730 ;
        RECT  0.475 2.070 3.060 2.730 ;
        RECT  0.305 1.800 0.475 2.730 ;
        RECT  0.000 2.070 0.305 2.730 ;
        END
    END VDD
END CELL104

MACRO CELL36
    CLASS CORE ;
    FOREIGN CELL36 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 2.400 ;
    SYMMETRY x y ;
    PIN QN
        ANTENNADIFFAREA 0.3444 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.670 0.710 5.750 1.490 ;
        RECT  5.650 0.495 5.670 1.905 ;
        RECT  5.560 0.495 5.650 0.890 ;
        RECT  5.560 1.310 5.650 1.905 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3360 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.150 0.790 5.195 0.900 ;
        RECT  5.045 0.790 5.150 1.490 ;
        RECT  4.985 0.790 5.045 0.900 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.1334 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.910 0.360 1.300 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0772 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.995 0.590 1.165 ;
        RECT  0.450 0.710 0.550 1.165 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0511 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 0.910 1.750 1.165 ;
        RECT  1.450 0.910 1.640 1.090 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.930 -0.330 6.000 0.330 ;
        RECT  5.820 -0.330 5.930 0.600 ;
        RECT  5.445 -0.330 5.820 0.330 ;
        RECT  5.255 -0.330 5.445 0.520 ;
        RECT  4.925 -0.330 5.255 0.330 ;
        RECT  4.735 -0.330 4.925 0.520 ;
        RECT  4.380 -0.330 4.735 0.330 ;
        RECT  4.190 -0.330 4.380 0.520 ;
        RECT  3.190 -0.330 4.190 0.330 ;
        RECT  3.080 -0.330 3.190 0.810 ;
        RECT  0.485 -0.330 3.080 0.330 ;
        RECT  0.315 -0.330 0.485 0.600 ;
        RECT  0.000 -0.330 0.315 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.930 2.070 6.000 2.730 ;
        RECT  5.820 1.600 5.930 2.730 ;
        RECT  5.405 2.070 5.820 2.730 ;
        RECT  5.295 1.800 5.405 2.730 ;
        RECT  4.885 2.070 5.295 2.730 ;
        RECT  4.775 1.800 4.885 2.730 ;
        RECT  4.380 2.070 4.775 2.730 ;
        RECT  4.190 1.890 4.380 2.730 ;
        RECT  3.210 2.070 4.190 2.730 ;
        RECT  3.040 1.800 3.210 2.730 ;
        RECT  0.475 2.070 3.040 2.730 ;
        RECT  0.305 1.800 0.475 2.730 ;
        RECT  0.000 2.070 0.305 2.730 ;
        END
    END VDD
END CELL36

MACRO CELL14
    CLASS CORE ;
    FOREIGN CELL14 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.400 ;
    SYMMETRY x y ;
    PIN QN
        ANTENNADIFFAREA 0.3360 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.070 0.710 6.150 1.490 ;
        RECT  6.050 0.495 6.070 1.900 ;
        RECT  5.960 0.495 6.050 0.890 ;
        RECT  5.960 1.310 6.050 1.900 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.3360 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.450 0.790 5.550 1.490 ;
        RECT  5.340 0.790 5.450 0.900 ;
        RECT  5.390 1.310 5.450 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.1600 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.180 1.290 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0613 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.755 1.180 0.970 1.290 ;
        RECT  0.650 1.180 0.755 1.690 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0512 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.040 0.910 2.150 1.165 ;
        RECT  1.850 0.910 2.040 1.090 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.1009 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 0.910 1.750 1.300 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.330 -0.330 6.400 0.330 ;
        RECT  6.220 -0.330 6.330 0.600 ;
        RECT  5.825 -0.330 6.220 0.330 ;
        RECT  5.635 -0.330 5.825 0.520 ;
        RECT  5.280 -0.330 5.635 0.330 ;
        RECT  5.090 -0.330 5.280 0.520 ;
        RECT  4.750 -0.330 5.090 0.330 ;
        RECT  4.560 -0.330 4.750 0.520 ;
        RECT  3.615 -0.330 4.560 0.330 ;
        RECT  3.505 -0.330 3.615 0.820 ;
        RECT  0.000 -0.330 3.505 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.330 2.070 6.400 2.730 ;
        RECT  6.220 1.600 6.330 2.730 ;
        RECT  5.825 2.070 6.220 2.730 ;
        RECT  5.635 1.860 5.825 2.730 ;
        RECT  5.280 2.070 5.635 2.730 ;
        RECT  5.090 1.860 5.280 2.730 ;
        RECT  4.735 2.070 5.090 2.730 ;
        RECT  4.545 1.860 4.735 2.730 ;
        RECT  3.615 2.070 4.545 2.730 ;
        RECT  3.445 1.800 3.615 2.730 ;
        RECT  0.455 2.070 3.445 2.730 ;
        RECT  0.345 1.800 0.455 2.730 ;
        RECT  0.000 2.070 0.345 2.730 ;
        END
    END VDD
END CELL14

MACRO CELL22
    CLASS CORE ;
    FOREIGN CELL22 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.400 BY 2.400 ;
    SYMMETRY x y ;
    PIN Q
        ANTENNADIFFAREA 0.2940 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.050 0.710 5.150 1.490 ;
        RECT  4.870 0.710 5.050 0.890 ;
        RECT  4.870 1.310 5.050 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.1334 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.910 0.360 1.300 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0772 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.995 0.590 1.165 ;
        RECT  0.450 0.710 0.550 1.165 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0511 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 0.910 1.750 1.165 ;
        RECT  1.450 0.910 1.640 1.090 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.240 -0.330 5.400 0.330 ;
        RECT  3.130 -0.330 3.240 0.810 ;
        RECT  0.485 -0.330 3.130 0.330 ;
        RECT  0.315 -0.330 0.485 0.600 ;
        RECT  0.000 -0.330 0.315 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.260 2.070 5.400 2.730 ;
        RECT  3.090 1.800 3.260 2.730 ;
        RECT  0.475 2.070 3.090 2.730 ;
        RECT  0.305 1.800 0.475 2.730 ;
        RECT  0.000 2.070 0.305 2.730 ;
        END
    END VDD
END CELL22

MACRO CELL74
    CLASS CORE ;
    FOREIGN CELL74 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 2.400 ;
    SYMMETRY x y ;
    PIN Q
        ANTENNADIFFAREA 0.3360 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.250 0.710 5.350 1.490 ;
        RECT  5.050 0.710 5.250 0.890 ;
        RECT  5.095 1.310 5.250 1.490 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.1334 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.910 0.360 1.300 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0772 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.995 0.590 1.165 ;
        RECT  0.450 0.710 0.550 1.165 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0511 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 0.910 1.750 1.165 ;
        RECT  1.450 0.910 1.640 1.090 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.260 -0.330 5.600 0.330 ;
        RECT  3.150 -0.330 3.260 0.810 ;
        RECT  0.485 -0.330 3.150 0.330 ;
        RECT  0.315 -0.330 0.485 0.600 ;
        RECT  0.000 -0.330 0.315 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.475 2.070 5.600 2.730 ;
        RECT  5.365 1.800 5.475 2.730 ;
        RECT  4.955 2.070 5.365 2.730 ;
        RECT  4.845 1.800 4.955 2.730 ;
        RECT  4.450 2.070 4.845 2.730 ;
        RECT  4.260 1.870 4.450 2.730 ;
        RECT  3.280 2.070 4.260 2.730 ;
        RECT  3.110 1.800 3.280 2.730 ;
        RECT  0.475 2.070 3.110 2.730 ;
        RECT  0.305 1.800 0.475 2.730 ;
        RECT  0.000 2.070 0.305 2.730 ;
        END
    END VDD
END CELL74

MACRO CELL9
    CLASS CORE ;
    FOREIGN CELL9 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.3248 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.710 1.350 1.690 ;
        RECT  1.000 0.710 1.250 0.800 ;
        RECT  1.235 1.510 1.250 1.690 ;
        RECT  1.050 1.510 1.235 1.890 ;
        RECT  0.890 0.430 1.000 0.800 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0960 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.910 1.150 1.290 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0514 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.910 0.570 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 0.910 0.350 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.255 -0.330 1.400 0.330 ;
        RECT  1.145 -0.330 1.255 0.600 ;
        RECT  0.735 -0.330 1.145 0.330 ;
        RECT  0.625 -0.330 0.735 0.600 ;
        RECT  0.215 -0.330 0.625 0.330 ;
        RECT  0.105 -0.330 0.215 0.600 ;
        RECT  0.000 -0.330 0.105 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.735 2.070 1.400 2.730 ;
        RECT  0.625 1.600 0.735 2.730 ;
        RECT  0.000 2.070 0.625 2.730 ;
        END
    END VDD
END CELL9

MACRO CELL59
    CLASS CORE ;
    FOREIGN CELL59 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.1626 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.510 1.150 1.490 ;
        RECT  0.950 0.510 1.050 0.690 ;
        RECT  0.795 1.400 1.050 1.490 ;
        RECT  0.690 1.400 0.795 1.800 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.780 0.910 0.950 1.290 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.910 0.380 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.535 -0.330 1.200 0.330 ;
        RECT  0.425 -0.330 0.535 0.600 ;
        RECT  0.000 -0.330 0.425 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.055 2.070 1.200 2.730 ;
        RECT  0.945 1.600 1.055 2.730 ;
        RECT  0.535 2.070 0.945 2.730 ;
        RECT  0.425 1.600 0.535 2.730 ;
        RECT  0.000 2.070 0.425 2.730 ;
        END
    END VDD
END CELL59

MACRO CELL1
    CLASS CORE ;
    FOREIGN CELL1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.3252 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.430 1.150 1.490 ;
        RECT  0.945 0.430 1.050 0.800 ;
        RECT  0.800 1.400 1.050 1.490 ;
        RECT  0.680 1.400 0.800 1.800 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.830 0.910 0.950 1.290 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0517 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.910 0.380 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.535 -0.330 1.200 0.330 ;
        RECT  0.425 -0.330 0.535 0.600 ;
        RECT  0.000 -0.330 0.425 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.055 2.070 1.200 2.730 ;
        RECT  0.945 1.600 1.055 2.730 ;
        RECT  0.535 2.070 0.945 2.730 ;
        RECT  0.425 1.600 0.535 2.730 ;
        RECT  0.000 2.070 0.425 2.730 ;
        END
    END VDD
END CELL1

MACRO CELL20
    CLASS CORE ;
    FOREIGN CELL20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.4881 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.430 1.350 1.800 ;
        RECT  1.190 0.430 1.250 0.800 ;
        RECT  1.190 1.400 1.250 1.800 ;
        RECT  0.770 1.400 1.190 1.500 ;
        RECT  0.650 1.400 0.770 1.800 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0978 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.910 1.160 1.290 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0978 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.830 0.910 0.950 1.290 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0491 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.205 0.910 0.350 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.495 -0.330 1.400 0.330 ;
        RECT  0.385 -0.330 0.495 0.600 ;
        RECT  0.000 -0.330 0.385 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.035 2.070 1.400 2.730 ;
        RECT  0.925 1.600 1.035 2.730 ;
        RECT  0.495 2.070 0.925 2.730 ;
        RECT  0.385 1.600 0.495 2.730 ;
        RECT  0.000 2.070 0.385 2.730 ;
        END
    END VDD
END CELL20

MACRO CELL93
    CLASS CORE ;
    FOREIGN CELL93 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.4872 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.510 1.550 1.690 ;
        RECT  1.415 0.510 1.450 0.890 ;
        RECT  0.595 1.600 1.450 1.690 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.0990 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 0.995 0.620 1.165 ;
        RECT  0.450 0.710 0.550 1.165 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0990 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.810 0.710 0.950 1.165 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0990 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.710 1.160 1.165 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0517 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.180 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.485 -0.330 1.600 0.330 ;
        RECT  0.375 -0.330 0.485 0.600 ;
        RECT  0.000 -0.330 0.375 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.525 2.070 1.600 2.730 ;
        RECT  1.415 1.800 1.525 2.730 ;
        RECT  1.005 2.070 1.415 2.730 ;
        RECT  0.895 1.800 1.005 2.730 ;
        RECT  0.485 2.070 0.895 2.730 ;
        RECT  0.375 1.600 0.485 2.730 ;
        RECT  0.000 2.070 0.375 2.730 ;
        END
    END VDD
END CELL93

MACRO CELL96
    CLASS CORE ;
    FOREIGN CELL96 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.3018 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.065 0.710 1.150 1.690 ;
        RECT  1.050 0.710 1.065 1.890 ;
        RECT  0.820 0.710 1.050 0.800 ;
        RECT  0.955 1.510 1.050 1.890 ;
        RECT  0.710 0.510 0.820 0.800 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.0792 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.815 0.910 0.950 1.290 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0509 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.910 0.380 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.080 -0.330 1.200 0.330 ;
        RECT  0.970 -0.330 1.080 0.600 ;
        RECT  0.535 -0.330 0.970 0.330 ;
        RECT  0.425 -0.330 0.535 0.600 ;
        RECT  0.000 -0.330 0.425 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.535 2.070 1.200 2.730 ;
        RECT  0.425 1.600 0.535 2.730 ;
        RECT  0.000 2.070 0.425 2.730 ;
        END
    END VDD
END CELL96

MACRO CELL5
    CLASS CORE ;
    FOREIGN CELL5 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.3228 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.255 0.710 1.350 1.690 ;
        RECT  1.250 0.710 1.255 1.890 ;
        RECT  1.245 0.710 1.250 0.800 ;
        RECT  1.155 1.510 1.250 1.890 ;
        RECT  1.135 0.510 1.245 0.800 ;
        RECT  0.750 0.710 1.135 0.800 ;
        RECT  0.620 0.510 0.750 0.800 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0792 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.005 0.910 1.155 1.290 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0792 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 1.000 0.835 1.170 ;
        RECT  0.650 1.000 0.750 1.290 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0508 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.200 0.910 0.350 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.015 -0.330 1.400 0.330 ;
        RECT  0.845 -0.330 1.015 0.600 ;
        RECT  0.495 -0.330 0.845 0.330 ;
        RECT  0.325 -0.330 0.495 0.600 ;
        RECT  0.000 -0.330 0.325 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.465 2.070 1.400 2.730 ;
        RECT  0.355 1.600 0.465 2.730 ;
        RECT  0.000 2.070 0.355 2.730 ;
        END
    END VDD
END CELL5

MACRO CELL86
    CLASS CORE ;
    FOREIGN CELL86 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.3078 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.505 0.710 1.550 1.690 ;
        RECT  1.450 0.710 1.505 1.890 ;
        RECT  1.260 0.710 1.450 0.800 ;
        RECT  1.395 1.510 1.450 1.890 ;
        RECT  1.150 0.510 1.260 0.800 ;
        RECT  0.750 0.710 1.150 0.800 ;
        RECT  0.640 0.510 0.750 0.800 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.0792 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 0.910 1.360 1.290 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0792 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.910 1.150 1.290 ;
        RECT  0.995 0.910 1.050 1.165 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0792 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.910 0.835 1.165 ;
        RECT  0.650 0.910 0.750 1.290 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.0508 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.190 0.910 0.350 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.520 -0.330 1.600 0.330 ;
        RECT  1.410 -0.330 1.520 0.600 ;
        RECT  1.000 -0.330 1.410 0.330 ;
        RECT  0.890 -0.330 1.000 0.600 ;
        RECT  0.465 -0.330 0.890 0.330 ;
        RECT  0.355 -0.330 0.465 0.600 ;
        RECT  0.000 -0.330 0.355 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.465 2.070 1.600 2.730 ;
        RECT  0.355 1.600 0.465 2.730 ;
        RECT  0.000 2.070 0.355 2.730 ;
        END
    END VDD
END CELL86

MACRO CELL41
    CLASS CORE ;
    FOREIGN CELL41 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.600 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.3408 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.510 0.550 1.890 ;
        RECT  0.380 0.510 0.450 0.890 ;
        RECT  0.380 1.310 0.450 1.890 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 1.000 0.245 1.170 ;
        RECT  0.050 1.000 0.150 1.290 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.225 -0.330 0.600 0.330 ;
        RECT  0.115 -0.330 0.225 0.800 ;
        RECT  0.000 -0.330 0.115 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.225 2.070 0.600 2.730 ;
        RECT  0.115 1.400 0.225 2.730 ;
        RECT  0.000 2.070 0.115 2.730 ;
        END
    END VDD
END CELL41

MACRO CELL35
    CLASS CORE ;
    FOREIGN CELL35 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.3360 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.455 0.710 0.550 1.490 ;
        RECT  0.450 0.510 0.455 1.890 ;
        RECT  0.345 0.510 0.450 0.890 ;
        RECT  0.345 1.310 0.450 1.890 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.2017 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.160 1.000 0.245 1.170 ;
        RECT  0.050 1.000 0.160 1.290 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.715 -0.330 0.800 0.330 ;
        RECT  0.605 -0.330 0.715 0.600 ;
        RECT  0.195 -0.330 0.605 0.330 ;
        RECT  0.085 -0.330 0.195 0.800 ;
        RECT  0.000 -0.330 0.085 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.715 2.070 0.800 2.730 ;
        RECT  0.605 1.600 0.715 2.730 ;
        RECT  0.195 2.070 0.605 2.730 ;
        RECT  0.085 1.400 0.195 2.730 ;
        RECT  0.000 2.070 0.085 2.730 ;
        END
    END VDD
END CELL35

MACRO CELL57
    CLASS CORE ;
    FOREIGN CELL57 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.3252 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.430 1.350 1.490 ;
        RECT  1.160 0.430 1.250 0.800 ;
        RECT  0.985 1.400 1.250 1.490 ;
        RECT  0.875 1.400 0.985 1.800 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.1009 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.910 1.160 1.290 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0514 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.910 0.555 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.910 0.350 1.290 ;
        RECT  0.180 1.000 0.250 1.170 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.725 -0.330 1.400 0.330 ;
        RECT  0.615 -0.330 0.725 0.600 ;
        RECT  0.000 -0.330 0.615 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.245 2.070 1.400 2.730 ;
        RECT  1.135 1.600 1.245 2.730 ;
        RECT  0.715 2.070 1.135 2.730 ;
        RECT  0.605 1.600 0.715 2.730 ;
        RECT  0.185 2.070 0.605 2.730 ;
        RECT  0.075 1.400 0.185 2.730 ;
        RECT  0.000 2.070 0.075 2.730 ;
        END
    END VDD
END CELL57

MACRO CELL112
    CLASS CORE ;
    FOREIGN CELL112 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.5280 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.460 1.310 1.575 1.890 ;
        RECT  1.450 0.710 1.460 1.890 ;
        RECT  1.360 0.710 1.450 1.690 ;
        RECT  1.130 0.710 1.360 0.800 ;
        RECT  1.055 1.510 1.360 1.690 ;
        RECT  0.945 1.510 1.055 1.890 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.2017 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.910 1.195 1.290 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.910 0.595 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.225 0.910 0.350 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.870 -0.330 2.000 0.330 ;
        RECT  1.760 -0.330 1.870 0.800 ;
        RECT  0.760 -0.330 1.760 0.330 ;
        RECT  0.650 -0.330 0.760 0.600 ;
        RECT  0.000 -0.330 0.650 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.845 2.070 2.000 2.730 ;
        RECT  1.735 1.400 1.845 2.730 ;
        RECT  1.315 2.070 1.735 2.730 ;
        RECT  1.205 1.800 1.315 2.730 ;
        RECT  0.795 2.070 1.205 2.730 ;
        RECT  0.685 1.600 0.795 2.730 ;
        RECT  0.240 2.070 0.685 2.730 ;
        RECT  0.130 1.400 0.240 2.730 ;
        RECT  0.000 2.070 0.130 2.730 ;
        END
    END VDD
END CELL112

MACRO CELL43
    CLASS CORE ;
    FOREIGN CELL43 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.3360 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.550 1.600 ;
        RECT  0.960 0.710 1.450 0.800 ;
        RECT  1.075 1.490 1.450 1.600 ;
        RECT  0.850 0.430 0.960 0.800 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.1009 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.910 0.560 1.300 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.180 1.290 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.1009 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 0.910 1.360 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1009 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.020 0.910 1.150 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.485 -0.330 1.600 0.330 ;
        RECT  1.375 -0.330 1.485 0.600 ;
        RECT  0.705 -0.330 1.375 0.330 ;
        RECT  0.595 -0.330 0.705 0.600 ;
        RECT  0.180 -0.330 0.595 0.330 ;
        RECT  0.070 -0.330 0.180 0.800 ;
        RECT  0.000 -0.330 0.070 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.705 2.070 1.600 2.730 ;
        RECT  0.595 1.400 0.705 2.730 ;
        RECT  0.000 2.070 0.595 2.730 ;
        END
    END VDD
END CELL43

MACRO CELL100
    CLASS CORE ;
    FOREIGN CELL100 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.3360 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.550 1.690 ;
        RECT  1.075 0.710 1.450 0.890 ;
        RECT  0.960 1.600 1.450 1.690 ;
        RECT  0.850 1.510 0.960 1.890 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.1009 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.900 0.560 1.290 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.180 1.290 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 1.000 1.360 1.490 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.000 1.150 1.490 ;
        RECT  1.020 1.000 1.050 1.170 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.705 -0.330 1.600 0.330 ;
        RECT  0.595 -0.330 0.705 0.780 ;
        RECT  0.000 -0.330 0.595 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.485 2.070 1.600 2.730 ;
        RECT  1.375 1.800 1.485 2.730 ;
        RECT  0.705 2.070 1.375 2.730 ;
        RECT  0.595 1.600 0.705 2.730 ;
        RECT  0.185 2.070 0.595 2.730 ;
        RECT  0.075 1.600 0.185 2.730 ;
        RECT  0.000 2.070 0.075 2.730 ;
        END
    END VDD
END CELL100

MACRO CELL94
    CLASS CORE ;
    FOREIGN CELL94 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 0.1344 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.620 0.510 1.750 1.910 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.1014 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 0.910 0.360 1.400 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.0507 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.210 0.710 1.350 1.290 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.0507 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.910 0.565 1.400 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.465 -0.330 1.800 0.330 ;
        RECT  1.355 -0.330 1.465 0.600 ;
        RECT  0.450 -0.330 1.355 0.330 ;
        RECT  0.340 -0.330 0.450 0.800 ;
        RECT  0.000 -0.330 0.340 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.465 2.070 1.800 2.730 ;
        RECT  1.355 1.800 1.465 2.730 ;
        RECT  0.450 2.070 1.355 2.730 ;
        RECT  0.340 1.800 0.450 2.730 ;
        RECT  0.000 2.070 0.340 2.730 ;
        END
    END VDD
END CELL94

MACRO CELL99
    CLASS CORE ;
    FOREIGN CELL99 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.1572 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.490 0.750 1.490 ;
        RECT  0.555 0.490 0.650 0.600 ;
        RECT  0.455 1.400 0.650 1.490 ;
        RECT  0.345 1.400 0.455 1.800 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.180 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.910 0.550 1.300 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.195 -0.330 0.800 0.330 ;
        RECT  0.085 -0.330 0.195 0.600 ;
        RECT  0.000 -0.330 0.085 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.715 2.070 0.800 2.730 ;
        RECT  0.605 1.600 0.715 2.730 ;
        RECT  0.195 2.070 0.605 2.730 ;
        RECT  0.085 1.400 0.195 2.730 ;
        RECT  0.000 2.070 0.085 2.730 ;
        END
    END VDD
END CELL99

MACRO CELL62
    CLASS CORE ;
    FOREIGN CELL62 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.3144 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.500 0.750 1.490 ;
        RECT  0.575 0.500 0.650 0.800 ;
        RECT  0.455 1.400 0.650 1.490 ;
        RECT  0.345 1.400 0.455 1.800 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.180 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.910 0.550 1.300 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.195 -0.330 0.800 0.330 ;
        RECT  0.085 -0.330 0.195 0.800 ;
        RECT  0.000 -0.330 0.085 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.715 2.070 0.800 2.730 ;
        RECT  0.605 1.600 0.715 2.730 ;
        RECT  0.195 2.070 0.605 2.730 ;
        RECT  0.085 1.600 0.195 2.730 ;
        RECT  0.000 2.070 0.085 2.730 ;
        END
    END VDD
END CELL62

MACRO CELL53
    CLASS CORE ;
    FOREIGN CELL53 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.5280 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 1.400 1.045 1.510 ;
        RECT  0.615 0.510 0.785 0.800 ;
        RECT  0.550 0.710 0.615 0.800 ;
        RECT  0.450 0.710 0.550 1.510 ;
        RECT  0.355 1.400 0.450 1.510 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.2016 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.220 1.000 1.350 1.690 ;
        RECT  0.180 1.600 1.220 1.690 ;
        RECT  0.050 1.000 0.180 1.690 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2017 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.910 0.760 1.300 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.275 -0.330 1.400 0.330 ;
        RECT  1.165 -0.330 1.275 0.800 ;
        RECT  0.235 -0.330 1.165 0.330 ;
        RECT  0.125 -0.330 0.235 0.800 ;
        RECT  0.000 -0.330 0.125 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.275 2.070 1.400 2.730 ;
        RECT  1.165 1.800 1.275 2.730 ;
        RECT  0.755 2.070 1.165 2.730 ;
        RECT  0.645 1.800 0.755 2.730 ;
        RECT  0.235 2.070 0.645 2.730 ;
        RECT  0.125 1.800 0.235 2.730 ;
        RECT  0.000 2.070 0.125 2.730 ;
        END
    END VDD
END CELL53

MACRO CELL15
    CLASS CORE ;
    FOREIGN CELL15 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.2682 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.490 1.150 1.490 ;
        RECT  0.850 0.490 1.050 0.600 ;
        RECT  0.935 1.400 1.050 1.800 ;
        RECT  0.550 1.400 0.935 1.490 ;
        RECT  0.420 1.400 0.550 1.800 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.230 0.910 0.350 1.290 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.910 0.605 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 0.910 0.950 1.300 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.270 -0.330 1.200 0.330 ;
        RECT  0.160 -0.330 0.270 0.600 ;
        RECT  0.000 -0.330 0.160 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.790 2.070 1.200 2.730 ;
        RECT  0.680 1.600 0.790 2.730 ;
        RECT  0.270 2.070 0.680 2.730 ;
        RECT  0.160 1.400 0.270 2.730 ;
        RECT  0.000 2.070 0.160 2.730 ;
        END
    END VDD
END CELL15

MACRO CELL105
    CLASS CORE ;
    FOREIGN CELL105 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.5364 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.510 1.150 1.490 ;
        RECT  0.895 0.510 1.050 0.800 ;
        RECT  1.035 1.400 1.050 1.490 ;
        RECT  0.920 1.400 1.035 1.800 ;
        RECT  0.550 1.400 0.920 1.490 ;
        RECT  0.390 1.400 0.550 1.800 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.910 0.360 1.290 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.910 0.590 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.825 0.910 0.950 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.255 -0.330 1.200 0.330 ;
        RECT  0.145 -0.330 0.255 0.800 ;
        RECT  0.000 -0.330 0.145 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.775 2.070 1.200 2.730 ;
        RECT  0.665 1.600 0.775 2.730 ;
        RECT  0.255 2.070 0.665 2.730 ;
        RECT  0.145 1.400 0.255 2.730 ;
        RECT  0.000 2.070 0.145 2.730 ;
        END
    END VDD
END CELL105

MACRO CELL90
    CLASS CORE ;
    FOREIGN CELL90 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.2640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.490 1.350 1.490 ;
        RECT  1.050 0.490 1.250 0.600 ;
        RECT  0.980 1.400 1.250 1.490 ;
        RECT  0.850 1.400 0.980 1.800 ;
        RECT  0.455 1.400 0.850 1.490 ;
        RECT  0.340 1.400 0.455 1.800 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.185 1.290 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.910 0.550 1.300 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.910 0.785 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.910 1.150 1.300 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.190 -0.330 1.400 0.330 ;
        RECT  0.080 -0.330 0.190 0.600 ;
        RECT  0.000 -0.330 0.080 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.230 2.070 1.400 2.730 ;
        RECT  1.120 1.600 1.230 2.730 ;
        RECT  0.710 2.070 1.120 2.730 ;
        RECT  0.600 1.600 0.710 2.730 ;
        RECT  0.190 2.070 0.600 2.730 ;
        RECT  0.080 1.400 0.190 2.730 ;
        RECT  0.000 2.070 0.080 2.730 ;
        END
    END VDD
END CELL90

MACRO CELL107
    CLASS CORE ;
    FOREIGN CELL107 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.5280 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.510 1.355 1.490 ;
        RECT  1.090 0.510 1.250 0.800 ;
        RECT  0.980 1.400 1.250 1.490 ;
        RECT  0.850 1.400 0.980 1.800 ;
        RECT  0.455 1.400 0.850 1.490 ;
        RECT  0.340 1.400 0.455 1.800 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.185 0.910 0.350 1.290 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.910 0.550 1.300 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.910 0.790 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.910 1.160 1.300 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.190 -0.330 1.400 0.330 ;
        RECT  0.080 -0.330 0.190 0.800 ;
        RECT  0.000 -0.330 0.080 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.230 2.070 1.400 2.730 ;
        RECT  1.120 1.600 1.230 2.730 ;
        RECT  0.710 2.070 1.120 2.730 ;
        RECT  0.600 1.600 0.710 2.730 ;
        RECT  0.190 2.070 0.600 2.730 ;
        RECT  0.080 1.400 0.190 2.730 ;
        RECT  0.000 2.070 0.080 2.730 ;
        END
    END VDD
END CELL107

MACRO CELL109
    CLASS CORE ;
    FOREIGN CELL109 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.1536 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.750 1.800 ;
        RECT  0.455 0.710 0.650 0.800 ;
        RECT  0.610 1.400 0.650 1.800 ;
        RECT  0.345 0.510 0.455 0.800 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.180 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.430 0.910 0.550 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.715 -0.330 0.800 0.330 ;
        RECT  0.605 -0.330 0.715 0.600 ;
        RECT  0.195 -0.330 0.605 0.330 ;
        RECT  0.085 -0.330 0.195 0.600 ;
        RECT  0.000 -0.330 0.085 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.195 2.070 0.800 2.730 ;
        RECT  0.085 1.400 0.195 2.730 ;
        RECT  0.000 2.070 0.085 2.730 ;
        END
    END VDD
END CELL109

MACRO CELL97
    CLASS CORE ;
    FOREIGN CELL97 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.3072 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.750 1.890 ;
        RECT  0.455 0.710 0.650 0.800 ;
        RECT  0.610 1.510 0.650 1.890 ;
        RECT  0.345 0.430 0.455 0.800 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.180 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.430 0.910 0.550 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.715 -0.330 0.800 0.330 ;
        RECT  0.605 -0.330 0.715 0.600 ;
        RECT  0.195 -0.330 0.605 0.330 ;
        RECT  0.085 -0.330 0.195 0.800 ;
        RECT  0.000 -0.330 0.085 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.195 2.070 0.800 2.730 ;
        RECT  0.085 1.600 0.195 2.730 ;
        RECT  0.000 2.070 0.085 2.730 ;
        END
    END VDD
END CELL97

MACRO CELL75
    CLASS CORE ;
    FOREIGN CELL75 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.4800 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.905 0.430 1.015 0.800 ;
        RECT  0.555 0.710 0.905 0.800 ;
        RECT  0.555 1.400 0.795 1.490 ;
        RECT  0.495 0.710 0.555 1.490 ;
        RECT  0.445 0.430 0.495 1.490 ;
        RECT  0.385 0.430 0.445 0.800 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.2018 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.135 0.910 1.155 1.490 ;
        RECT  1.045 0.910 1.135 1.690 ;
        RECT  0.355 1.600 1.045 1.690 ;
        RECT  0.265 0.910 0.355 1.690 ;
        RECT  0.245 0.910 0.265 1.490 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2017 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.645 0.910 0.760 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.275 -0.330 1.400 0.330 ;
        RECT  1.165 -0.330 1.275 0.800 ;
        RECT  0.765 -0.330 1.165 0.330 ;
        RECT  0.635 -0.330 0.765 0.600 ;
        RECT  0.235 -0.330 0.635 0.330 ;
        RECT  0.125 -0.330 0.235 0.800 ;
        RECT  0.000 -0.330 0.125 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.335 2.070 1.400 2.730 ;
        RECT  1.225 1.600 1.335 2.730 ;
        RECT  0.175 2.070 1.225 2.730 ;
        RECT  0.075 1.600 0.175 2.730 ;
        RECT  0.000 2.070 0.075 2.730 ;
        END
    END VDD
END CELL75

MACRO CELL33
    CLASS CORE ;
    FOREIGN CELL33 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.2352 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.710 0.750 1.890 ;
        RECT  0.455 0.710 0.650 0.800 ;
        RECT  0.610 1.510 0.650 1.890 ;
        RECT  0.345 0.510 0.455 0.800 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.0792 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.180 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0792 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.430 0.910 0.550 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.715 -0.330 0.800 0.330 ;
        RECT  0.605 -0.330 0.715 0.600 ;
        RECT  0.195 -0.330 0.605 0.330 ;
        RECT  0.085 -0.330 0.195 0.600 ;
        RECT  0.000 -0.330 0.085 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.195 2.070 0.800 2.730 ;
        RECT  0.085 1.600 0.195 2.730 ;
        RECT  0.000 2.070 0.085 2.730 ;
        END
    END VDD
END CELL33

MACRO CELL12
    CLASS CORE ;
    FOREIGN CELL12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.3426 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.710 1.150 1.690 ;
        RECT  1.035 0.710 1.045 0.800 ;
        RECT  1.035 1.510 1.045 1.690 ;
        RECT  0.925 0.510 1.035 0.800 ;
        RECT  0.850 1.510 1.035 1.890 ;
        RECT  0.515 0.710 0.925 0.800 ;
        RECT  0.405 0.510 0.515 0.800 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.0792 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.350 1.090 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0792 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.910 0.600 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0792 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.830 0.910 0.950 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.775 -0.330 1.200 0.330 ;
        RECT  0.665 -0.330 0.775 0.600 ;
        RECT  0.255 -0.330 0.665 0.330 ;
        RECT  0.145 -0.330 0.255 0.600 ;
        RECT  0.000 -0.330 0.145 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.255 2.070 1.200 2.730 ;
        RECT  0.145 1.400 0.255 2.730 ;
        RECT  0.000 2.070 0.145 2.730 ;
        END
    END VDD
END CELL12

MACRO CELL32
    CLASS CORE ;
    FOREIGN CELL32 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.3360 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.710 1.350 1.690 ;
        RECT  0.975 0.710 1.250 0.800 ;
        RECT  1.235 1.510 1.250 1.690 ;
        RECT  1.050 1.510 1.235 1.890 ;
        RECT  0.865 0.510 0.975 0.800 ;
        RECT  0.455 0.710 0.865 0.800 ;
        RECT  0.345 0.510 0.455 0.800 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.0792 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.350 1.090 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0792 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.910 0.555 1.290 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0792 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.910 0.790 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0792 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.910 1.160 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.235 -0.330 1.400 0.330 ;
        RECT  1.125 -0.330 1.235 0.600 ;
        RECT  0.715 -0.330 1.125 0.330 ;
        RECT  0.605 -0.330 0.715 0.600 ;
        RECT  0.195 -0.330 0.605 0.330 ;
        RECT  0.085 -0.330 0.195 0.600 ;
        RECT  0.000 -0.330 0.085 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.195 2.070 1.400 2.730 ;
        RECT  0.085 1.400 0.195 2.730 ;
        RECT  0.000 2.070 0.085 2.730 ;
        END
    END VDD
END CELL32

MACRO CELL54
    CLASS CORE ;
    FOREIGN CELL54 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 0.3360 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.490 1.550 1.710 ;
        RECT  1.345 0.490 1.450 0.590 ;
        RECT  1.335 1.600 1.450 1.710 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.020 0.910 1.150 1.290 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.910 0.785 1.290 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.180 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.910 0.550 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.225 -0.330 1.600 0.330 ;
        RECT  1.115 -0.330 1.225 0.590 ;
        RECT  0.000 -0.330 1.115 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.225 2.070 1.600 2.730 ;
        RECT  1.115 1.600 1.225 2.730 ;
        RECT  0.705 2.070 1.115 2.730 ;
        RECT  0.595 1.600 0.705 2.730 ;
        RECT  0.000 2.070 0.595 2.730 ;
        END
    END VDD
END CELL54

MACRO CELL58
    CLASS CORE ;
    FOREIGN CELL58 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 0.4200 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.260 0.710 1.350 1.490 ;
        RECT  1.250 0.510 1.260 1.890 ;
        RECT  1.145 0.510 1.250 0.890 ;
        RECT  1.145 1.310 1.250 1.890 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.910 0.800 1.290 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.170 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.430 0.910 0.550 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.975 -0.330 1.400 0.330 ;
        RECT  0.865 -0.330 0.975 0.600 ;
        RECT  0.000 -0.330 0.865 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.975 2.070 1.400 2.730 ;
        RECT  0.865 1.600 0.975 2.730 ;
        RECT  0.195 2.070 0.865 2.730 ;
        RECT  0.085 1.600 0.195 2.730 ;
        RECT  0.000 2.070 0.085 2.730 ;
        END
    END VDD
END CELL58

MACRO CELL80
    CLASS CORE ;
    FOREIGN CELL80 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 0.2688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.510 1.950 1.940 ;
        RECT  1.820 0.510 1.850 0.890 ;
        RECT  1.780 1.800 1.850 1.940 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.415 1.000 1.550 1.490 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 1.000 1.235 1.170 ;
        RECT  1.050 1.000 1.150 1.490 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 1.000 0.960 1.490 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.170 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 1.000 0.550 1.490 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.670 -0.330 2.000 0.330 ;
        RECT  1.560 -0.330 1.670 0.800 ;
        RECT  0.000 -0.330 1.560 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.670 2.070 2.000 2.730 ;
        RECT  1.560 1.800 1.670 2.730 ;
        RECT  0.170 2.070 1.560 2.730 ;
        RECT  0.060 1.600 0.170 2.730 ;
        RECT  0.000 2.070 0.060 2.730 ;
        END
    END VDD
END CELL80

MACRO CELL29
    CLASS CORE ;
    FOREIGN CELL29 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 0.2688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.625 0.510 1.750 1.890 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.910 0.560 1.290 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.180 1.290 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.910 0.770 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.035 0.910 1.150 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.470 -0.330 1.800 0.330 ;
        RECT  1.360 -0.330 1.470 0.600 ;
        RECT  0.440 -0.330 1.360 0.330 ;
        RECT  0.330 -0.330 0.440 0.590 ;
        RECT  0.000 -0.330 0.330 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.475 2.070 1.800 2.730 ;
        RECT  1.355 1.600 1.475 2.730 ;
        RECT  0.705 2.070 1.355 2.730 ;
        RECT  0.585 1.600 0.705 2.730 ;
        RECT  0.000 2.070 0.585 2.730 ;
        END
    END VDD
END CELL29

MACRO CELL66
    CLASS CORE ;
    FOREIGN CELL66 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 0.3360 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.510 1.550 1.890 ;
        RECT  1.375 0.510 1.450 0.890 ;
        RECT  1.375 1.710 1.450 1.890 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.910 1.150 1.290 ;
        RECT  0.920 1.025 1.040 1.135 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.910 0.790 1.290 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.910 0.560 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.170 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.225 -0.330 1.600 0.330 ;
        RECT  1.115 -0.330 1.225 0.800 ;
        RECT  0.000 -0.330 1.115 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.225 2.070 1.600 2.730 ;
        RECT  1.115 1.600 1.225 2.730 ;
        RECT  0.185 2.070 1.115 2.730 ;
        RECT  0.075 1.600 0.185 2.730 ;
        RECT  0.000 2.070 0.075 2.730 ;
        END
    END VDD
END CELL66

MACRO CELL7
    CLASS CORE ;
    FOREIGN CELL7 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 0.1470 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.490 1.950 1.890 ;
        RECT  1.760 0.490 1.850 0.600 ;
        RECT  1.810 1.710 1.850 1.890 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.910 0.550 1.290 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.170 1.290 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0509 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 1.110 0.770 1.490 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0512 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.025 1.110 1.150 1.490 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0508 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.245 1.110 1.360 1.490 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.650 -0.330 2.000 0.330 ;
        RECT  1.540 -0.330 1.650 0.600 ;
        RECT  0.445 -0.330 1.540 0.330 ;
        RECT  0.335 -0.330 0.445 0.600 ;
        RECT  0.000 -0.330 0.335 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.560 2.070 2.000 2.730 ;
        RECT  1.450 1.800 1.560 2.730 ;
        RECT  0.185 2.070 1.450 2.730 ;
        RECT  0.075 1.600 0.185 2.730 ;
        RECT  0.000 2.070 0.075 2.730 ;
        END
    END VDD
END CELL7

MACRO CELL37
    CLASS CORE ;
    FOREIGN CELL37 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 0.2688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.820 0.510 1.950 1.890 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.035 0.910 1.150 1.290 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.910 1.385 1.290 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.910 0.790 1.290 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.910 0.560 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.170 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.220 -0.330 2.000 0.330 ;
        RECT  1.120 -0.330 1.220 0.600 ;
        RECT  0.000 -0.330 1.120 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.575 2.070 2.000 2.730 ;
        RECT  1.465 1.600 1.575 2.730 ;
        RECT  0.185 2.070 1.465 2.730 ;
        RECT  0.075 1.600 0.185 2.730 ;
        RECT  0.000 2.070 0.075 2.730 ;
        END
    END VDD
END CELL37

MACRO CELL92
    CLASS CORE ;
    FOREIGN CELL92 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.4992 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.690 1.350 1.490 ;
        RECT  0.305 0.690 1.250 0.780 ;
        RECT  0.970 1.400 1.250 1.490 ;
        RECT  0.850 1.400 0.970 1.800 ;
        RECT  0.190 1.400 0.850 1.490 ;
        RECT  0.050 1.400 0.190 1.800 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.910 1.160 1.290 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.910 0.790 1.290 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.170 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.910 0.560 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.235 -0.330 1.400 0.330 ;
        RECT  1.125 -0.330 1.235 0.600 ;
        RECT  0.000 -0.330 1.125 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.235 2.070 1.400 2.730 ;
        RECT  1.125 1.600 1.235 2.730 ;
        RECT  0.715 2.070 1.125 2.730 ;
        RECT  0.605 1.600 0.715 2.730 ;
        RECT  0.000 2.070 0.605 2.730 ;
        END
    END VDD
END CELL92

MACRO CELL8
    CLASS CORE ;
    FOREIGN CELL8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.1860 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.685 1.150 1.490 ;
        RECT  0.375 0.685 1.050 0.775 ;
        RECT  0.770 1.400 1.050 1.490 ;
        RECT  0.650 1.400 0.770 1.800 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.805 0.910 0.950 1.290 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.220 0.910 0.350 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.910 0.585 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.085 -0.330 1.200 0.330 ;
        RECT  0.975 -0.330 1.085 0.595 ;
        RECT  0.000 -0.330 0.975 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.030 2.070 1.200 2.730 ;
        RECT  0.920 1.600 1.030 2.730 ;
        RECT  0.255 2.070 0.920 2.730 ;
        RECT  0.135 1.400 0.255 2.730 ;
        RECT  0.000 2.070 0.135 2.730 ;
        END
    END VDD
END CELL8

MACRO CELL50
    CLASS CORE ;
    FOREIGN CELL50 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.3360 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.690 1.150 1.500 ;
        RECT  0.365 0.690 1.050 0.780 ;
        RECT  0.765 1.400 1.050 1.500 ;
        RECT  0.650 1.400 0.765 1.800 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.830 0.910 0.950 1.290 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.230 0.910 0.350 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.910 0.590 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.035 -0.330 1.200 0.330 ;
        RECT  0.925 -0.330 1.035 0.590 ;
        RECT  0.000 -0.330 0.925 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.035 2.070 1.200 2.730 ;
        RECT  0.925 1.600 1.035 2.730 ;
        RECT  0.260 2.070 0.925 2.730 ;
        RECT  0.140 1.400 0.260 2.730 ;
        RECT  0.000 2.070 0.140 2.730 ;
        END
    END VDD
END CELL50

MACRO CELL72
    CLASS CORE ;
    FOREIGN CELL72 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.2448 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.430 1.670 1.550 1.890 ;
        RECT  0.150 1.670 1.430 1.760 ;
        RECT  0.150 0.680 0.995 0.770 ;
        RECT  0.050 0.680 0.150 1.760 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.890 0.360 1.290 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.0513 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 1.110 0.565 1.490 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0513 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.440 0.800 1.550 1.560 ;
        RECT  0.840 1.470 1.440 1.560 ;
        RECT  0.655 1.400 0.840 1.560 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0511 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.020 0.910 1.150 1.380 ;
        RECT  0.655 0.910 1.020 1.060 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0509 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 0.800 1.350 1.330 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.180 -0.330 1.600 0.330 ;
        RECT  0.070 -0.330 0.180 0.590 ;
        RECT  0.000 -0.330 0.070 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.990 2.070 1.600 2.730 ;
        RECT  0.880 1.870 0.990 2.730 ;
        RECT  0.185 2.070 0.880 2.730 ;
        RECT  0.075 1.870 0.185 2.730 ;
        RECT  0.000 2.070 0.075 2.730 ;
        END
    END VDD
END CELL72

MACRO CELL65
    CLASS CORE ;
    FOREIGN CELL65 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.800 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.2448 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.620 1.670 1.750 1.890 ;
        RECT  0.350 1.670 1.620 1.770 ;
        RECT  0.865 0.680 1.245 0.770 ;
        RECT  0.775 0.680 0.865 0.890 ;
        RECT  0.350 0.800 0.775 0.890 ;
        RECT  0.250 0.800 0.350 1.770 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 1.100 0.560 1.490 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.900 0.160 1.290 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.0513 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.755 1.055 0.835 1.225 ;
        RECT  0.650 1.055 0.755 1.490 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0512 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 0.800 1.750 1.560 ;
        RECT  1.065 1.470 1.640 1.560 ;
        RECT  0.955 1.285 1.065 1.560 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.0510 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.210 0.910 1.350 1.380 ;
        RECT  1.030 0.910 1.210 1.090 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0509 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.440 0.910 1.550 1.330 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.485 -0.330 1.800 0.330 ;
        RECT  0.310 -0.330 0.485 0.530 ;
        RECT  0.000 -0.330 0.310 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.200 2.070 1.800 2.730 ;
        RECT  1.090 1.880 1.200 2.730 ;
        RECT  0.180 2.070 1.090 2.730 ;
        RECT  0.070 1.880 0.180 2.730 ;
        RECT  0.000 2.070 0.070 2.730 ;
        END
    END VDD
END CELL65

MACRO CELL40
    CLASS CORE ;
    FOREIGN CELL40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.5088 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.680 1.350 1.490 ;
        RECT  0.830 0.680 1.250 0.780 ;
        RECT  1.240 1.400 1.250 1.490 ;
        RECT  1.130 1.400 1.240 1.800 ;
        RECT  0.190 1.400 1.130 1.490 ;
        RECT  0.050 1.400 0.190 1.800 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.910 0.560 1.290 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.170 1.290 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.910 0.795 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.910 1.155 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.460 -0.330 1.400 0.330 ;
        RECT  0.350 -0.330 0.460 0.600 ;
        RECT  0.000 -0.330 0.350 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.720 2.070 1.400 2.730 ;
        RECT  0.610 1.600 0.720 2.730 ;
        RECT  0.000 2.070 0.610 2.730 ;
        END
    END VDD
END CELL40

MACRO CELL10
    CLASS CORE ;
    FOREIGN CELL10 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.6720 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 0.680 2.350 1.490 ;
        RECT  1.340 0.680 2.250 0.770 ;
        RECT  1.750 1.400 2.250 1.490 ;
        RECT  1.640 1.400 1.750 1.800 ;
        RECT  0.750 1.400 1.640 1.490 ;
        RECT  0.610 1.400 0.750 1.800 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.2017 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.910 1.150 1.310 ;
        RECT  0.170 1.220 1.030 1.310 ;
        RECT  0.050 0.910 0.170 1.310 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2017 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.910 0.750 1.130 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.2017 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 0.910 2.150 1.310 ;
        RECT  1.370 1.220 2.050 1.310 ;
        RECT  1.250 0.910 1.370 1.310 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2017 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.910 1.950 1.130 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.970 -0.330 2.400 0.330 ;
        RECT  0.860 -0.330 0.970 0.600 ;
        RECT  0.450 -0.330 0.860 0.330 ;
        RECT  0.340 -0.330 0.450 0.600 ;
        RECT  0.000 -0.330 0.340 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.270 2.070 2.400 2.730 ;
        RECT  2.160 1.600 2.270 2.730 ;
        RECT  1.230 2.070 2.160 2.730 ;
        RECT  1.120 1.600 1.230 2.730 ;
        RECT  0.190 2.070 1.120 2.730 ;
        RECT  0.080 1.600 0.190 2.730 ;
        RECT  0.000 2.070 0.080 2.730 ;
        END
    END VDD
END CELL10

MACRO CELL46
    CLASS CORE ;
    FOREIGN CELL46 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 1.4090 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.355 1.300 4.465 1.690 ;
        RECT  3.945 1.300 4.355 1.400 ;
        RECT  3.835 1.300 3.945 1.690 ;
        RECT  2.260 1.300 3.835 1.400 ;
        RECT  2.150 0.690 2.260 1.400 ;
        RECT  0.850 0.690 2.150 0.800 ;
        RECT  0.850 1.310 0.965 1.690 ;
        RECT  0.550 0.690 0.850 1.470 ;
        RECT  0.045 0.690 0.550 0.800 ;
        RECT  0.450 1.310 0.550 1.470 ;
        RECT  0.335 1.310 0.450 1.690 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.4034 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.970 3.150 1.130 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4034 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.850 0.970 4.350 1.130 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.4034 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.970 1.950 1.130 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4034 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.385 1.130 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.725 -0.330 4.800 0.330 ;
        RECT  4.615 -0.330 4.725 0.800 ;
        RECT  4.205 -0.330 4.615 0.330 ;
        RECT  4.095 -0.330 4.205 0.600 ;
        RECT  3.235 -0.330 4.095 0.330 ;
        RECT  3.125 -0.330 3.235 0.600 ;
        RECT  2.715 -0.330 3.125 0.330 ;
        RECT  2.605 -0.330 2.715 0.600 ;
        RECT  0.000 -0.330 2.605 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.975 2.070 4.800 2.730 ;
        RECT  2.865 1.800 2.975 2.730 ;
        RECT  2.455 2.070 2.865 2.730 ;
        RECT  2.345 1.600 2.455 2.730 ;
        RECT  1.935 2.070 2.345 2.730 ;
        RECT  1.825 1.800 1.935 2.730 ;
        RECT  0.000 2.070 1.825 2.730 ;
        END
    END VDD
END CELL46

MACRO CELL56
    CLASS CORE ;
    FOREIGN CELL56 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.4512 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.680 1.350 1.490 ;
        RECT  0.210 0.680 1.250 0.775 ;
        RECT  0.980 1.400 1.250 1.490 ;
        RECT  0.850 1.400 0.980 1.800 ;
        RECT  0.050 0.510 0.210 0.775 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.025 0.910 1.150 1.290 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.910 0.805 1.290 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.910 0.560 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.180 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.250 -0.330 1.400 0.330 ;
        RECT  1.140 -0.330 1.250 0.590 ;
        RECT  0.000 -0.330 1.140 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.250 2.070 1.400 2.730 ;
        RECT  1.140 1.600 1.250 2.730 ;
        RECT  0.210 2.070 1.140 2.730 ;
        RECT  0.100 1.600 0.210 2.730 ;
        RECT  0.000 2.070 0.100 2.730 ;
        END
    END VDD
END CELL56

MACRO CELL111
    CLASS CORE ;
    FOREIGN CELL111 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.600 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 1.6970 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.160 1.300 4.270 1.890 ;
        RECT  3.750 1.300 4.160 1.400 ;
        RECT  3.640 1.000 3.750 1.890 ;
        RECT  3.310 1.000 3.640 1.110 ;
        RECT  3.200 0.690 3.310 1.110 ;
        RECT  0.850 0.690 3.200 0.800 ;
        RECT  0.850 1.310 0.960 1.690 ;
        RECT  0.550 0.690 0.850 1.490 ;
        RECT  0.180 0.690 0.550 0.800 ;
        RECT  0.450 1.310 0.550 1.490 ;
        RECT  0.330 1.310 0.450 1.690 ;
        RECT  0.070 0.510 0.180 0.800 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.4034 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.995 0.910 4.405 1.130 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.4034 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.405 1.130 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4034 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.595 0.910 2.005 1.130 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4034 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.595 0.910 3.005 1.130 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.270 -0.330 4.600 0.330 ;
        RECT  4.160 -0.330 4.270 0.600 ;
        RECT  3.750 -0.330 4.160 0.330 ;
        RECT  3.640 -0.330 3.750 0.600 ;
        RECT  0.000 -0.330 3.640 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.530 2.070 4.600 2.730 ;
        RECT  4.420 1.400 4.530 2.730 ;
        RECT  4.010 2.070 4.420 2.730 ;
        RECT  3.900 1.600 4.010 2.730 ;
        RECT  3.490 2.070 3.900 2.730 ;
        RECT  3.380 1.400 3.490 2.730 ;
        RECT  2.970 2.070 3.380 2.730 ;
        RECT  2.860 1.600 2.970 2.730 ;
        RECT  0.000 2.070 2.860 2.730 ;
        END
    END VDD
END CELL111

MACRO CELL25
    CLASS CORE ;
    FOREIGN CELL25 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.2346 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 1.400 0.970 1.890 ;
        RECT  0.150 1.400 0.850 1.490 ;
        RECT  0.170 0.690 0.765 0.780 ;
        RECT  0.150 0.510 0.170 0.780 ;
        RECT  0.050 0.510 0.150 1.490 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.910 1.160 1.290 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.910 1.385 1.290 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.790 0.910 0.950 1.290 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.910 0.580 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.910 0.360 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.270 -0.330 1.600 0.330 ;
        RECT  1.160 -0.330 1.270 0.600 ;
        RECT  0.000 -0.330 1.160 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.500 2.070 1.600 2.730 ;
        RECT  1.390 1.600 1.500 2.730 ;
        RECT  0.200 2.070 1.390 2.730 ;
        RECT  0.090 1.600 0.200 2.730 ;
        RECT  0.000 2.070 0.090 2.730 ;
        END
    END VDD
END CELL25

MACRO CELL18
    CLASS CORE ;
    FOREIGN CELL18 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.4548 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 1.400 0.970 1.800 ;
        RECT  0.150 1.400 0.850 1.490 ;
        RECT  0.190 0.680 0.750 0.770 ;
        RECT  0.150 0.510 0.190 0.770 ;
        RECT  0.050 0.510 0.150 1.490 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.910 1.160 1.290 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.910 1.385 1.290 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.795 0.910 0.950 1.290 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1009 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.910 0.580 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1009 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.910 0.360 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.230 -0.330 1.600 0.330 ;
        RECT  1.120 -0.330 1.230 0.590 ;
        RECT  0.000 -0.330 1.120 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.490 2.070 1.600 2.730 ;
        RECT  1.380 1.400 1.490 2.730 ;
        RECT  0.190 2.070 1.380 2.730 ;
        RECT  0.080 1.600 0.190 2.730 ;
        RECT  0.000 2.070 0.080 2.730 ;
        END
    END VDD
END CELL18

MACRO CELL30
    CLASS CORE ;
    FOREIGN CELL30 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.2418 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 1.400 1.055 1.690 ;
        RECT  0.350 1.400 0.945 1.490 ;
        RECT  0.350 0.680 0.835 0.780 ;
        RECT  0.270 0.680 0.350 1.490 ;
        RECT  0.250 0.510 0.270 1.490 ;
        RECT  0.160 0.510 0.250 0.780 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.910 1.160 1.290 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.910 1.390 1.290 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.635 0.910 1.750 1.290 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.800 0.910 0.950 1.290 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.910 0.600 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0504 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.890 0.160 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.835 -0.330 2.000 0.330 ;
        RECT  1.725 -0.330 1.835 0.705 ;
        RECT  1.315 -0.330 1.725 0.330 ;
        RECT  1.205 -0.330 1.315 0.600 ;
        RECT  0.000 -0.330 1.205 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.835 2.070 2.000 2.730 ;
        RECT  1.725 1.400 1.835 2.730 ;
        RECT  0.275 2.070 1.725 2.730 ;
        RECT  0.165 1.600 0.275 2.730 ;
        RECT  0.000 2.070 0.165 2.730 ;
        END
    END VDD
END CELL30

MACRO CELL52
    CLASS CORE ;
    FOREIGN CELL52 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.4836 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.945 1.400 1.055 1.800 ;
        RECT  0.350 1.400 0.945 1.490 ;
        RECT  0.350 0.690 0.840 0.780 ;
        RECT  0.270 0.690 0.350 1.490 ;
        RECT  0.250 0.510 0.270 1.490 ;
        RECT  0.165 0.510 0.250 0.780 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.910 1.160 1.290 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 0.910 1.390 1.290 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 0.910 1.755 1.290 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.1009 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.800 0.910 0.950 1.290 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.910 0.610 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.890 0.160 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.835 -0.330 2.000 0.330 ;
        RECT  1.720 -0.330 1.835 0.780 ;
        RECT  1.315 -0.330 1.720 0.330 ;
        RECT  1.205 -0.330 1.315 0.600 ;
        RECT  0.000 -0.330 1.205 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.835 2.070 2.000 2.730 ;
        RECT  1.725 1.400 1.835 2.730 ;
        RECT  0.275 2.070 1.725 2.730 ;
        RECT  0.165 1.600 0.275 2.730 ;
        RECT  0.000 2.070 0.165 2.730 ;
        END
    END VDD
END CELL52

MACRO CELL88
    CLASS CORE ;
    FOREIGN CELL88 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 0.3444 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.055 0.710 1.150 1.490 ;
        RECT  1.050 0.510 1.055 1.890 ;
        RECT  0.945 0.510 1.050 0.890 ;
        RECT  0.945 1.310 1.050 1.890 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.0800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.910 0.610 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0792 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.910 0.360 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.795 -0.330 1.200 0.330 ;
        RECT  0.685 -0.330 0.795 0.600 ;
        RECT  0.250 -0.330 0.685 0.330 ;
        RECT  0.140 -0.330 0.250 0.800 ;
        RECT  0.000 -0.330 0.140 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.795 2.070 1.200 2.730 ;
        RECT  0.685 1.600 0.795 2.730 ;
        RECT  0.000 2.070 0.685 2.730 ;
        END
    END VDD
END CELL88

MACRO CELL102
    CLASS CORE ;
    FOREIGN CELL102 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 0.3108 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.490 1.550 1.890 ;
        RECT  1.350 0.490 1.450 0.600 ;
        RECT  1.420 1.310 1.450 1.890 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.0792 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.180 1.290 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.0792 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.435 0.910 0.560 1.290 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.0792 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 0.910 0.785 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.0800 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.020 0.910 1.150 1.290 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.240 -0.330 1.600 0.330 ;
        RECT  1.130 -0.330 1.240 0.600 ;
        RECT  0.720 -0.330 1.130 0.330 ;
        RECT  0.610 -0.330 0.720 0.600 ;
        RECT  0.200 -0.330 0.610 0.330 ;
        RECT  0.090 -0.330 0.200 0.600 ;
        RECT  0.000 -0.330 0.090 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.240 2.070 1.600 2.730 ;
        RECT  1.130 1.600 1.240 2.730 ;
        RECT  0.000 2.070 1.130 2.730 ;
        END
    END VDD
END CELL102

MACRO CELL27
    CLASS CORE ;
    FOREIGN CELL27 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.600 BY 2.400 ;
    SYMMETRY x y ;
    PIN SI
        ANTENNAGATEAREA 0.0188 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.560 1.100 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.0866 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.890 2.950 1.290 ;
        RECT  2.615 0.890 2.850 1.000 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.2688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.420 0.510 6.550 1.890 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.180 1.290 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.0505 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.790 0.810 0.900 ;
        RECT  0.635 0.510 0.750 0.900 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.0512 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.280 0.910 3.390 1.165 ;
        RECT  3.050 0.910 3.280 1.090 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.270 -0.330 6.600 0.330 ;
        RECT  6.160 -0.330 6.270 0.600 ;
        RECT  5.830 -0.330 6.160 0.330 ;
        RECT  5.660 -0.330 5.830 0.380 ;
        RECT  2.210 -0.330 5.660 0.330 ;
        RECT  2.100 -0.330 2.210 0.570 ;
        RECT  1.460 -0.330 2.100 0.330 ;
        RECT  1.290 -0.330 1.460 0.380 ;
        RECT  0.440 -0.330 1.290 0.330 ;
        RECT  0.330 -0.330 0.440 0.600 ;
        RECT  0.000 -0.330 0.330 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.270 2.070 6.600 2.730 ;
        RECT  6.160 1.790 6.270 2.730 ;
        RECT  4.835 2.070 6.160 2.730 ;
        RECT  4.665 1.800 4.835 2.730 ;
        RECT  0.440 2.070 4.665 2.730 ;
        RECT  0.330 1.600 0.440 2.730 ;
        RECT  0.000 2.070 0.330 2.730 ;
        END
    END VDD
END CELL27

MACRO CELL110
    CLASS CORE ;
    FOREIGN CELL110 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.600 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 0.1920 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 1.110 0.550 1.890 ;
        RECT  0.410 1.310 0.450 1.890 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.225 -0.330 0.600 0.330 ;
        RECT  0.115 -0.330 0.225 0.600 ;
        RECT  0.000 -0.330 0.115 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.225 2.070 0.600 2.730 ;
        RECT  0.115 1.400 0.225 2.730 ;
        RECT  0.000 2.070 0.115 2.730 ;
        END
    END VDD
END CELL110

MACRO CELL44
    CLASS CORE ;
    FOREIGN CELL44 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.600 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.1440 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 0.510 0.550 1.090 ;
        RECT  0.380 0.510 0.450 0.890 ;
        END
    END ZN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.225 -0.330 0.600 0.330 ;
        RECT  0.115 -0.330 0.225 0.800 ;
        RECT  0.000 -0.330 0.115 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.225 2.070 0.600 2.730 ;
        RECT  0.115 1.400 0.225 2.730 ;
        RECT  0.000 2.070 0.115 2.730 ;
        END
    END VDD
END CELL44

MACRO CELL108
    CLASS CORE ;
    FOREIGN CELL108 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.2940 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 0.710 1.950 1.690 ;
        RECT  1.850 0.710 1.855 1.890 ;
        RECT  1.830 0.710 1.850 0.890 ;
        RECT  1.745 1.510 1.850 1.890 ;
        RECT  1.720 0.510 1.830 0.890 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.1009 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.550 1.150 ;
        RECT  1.325 0.980 1.450 1.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1106 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.995 0.365 1.490 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.565 -0.330 2.000 0.330 ;
        RECT  1.435 -0.330 1.565 0.600 ;
        RECT  0.360 -0.330 1.435 0.330 ;
        RECT  0.360 0.745 0.475 0.855 ;
        RECT  0.270 -0.330 0.360 0.855 ;
        RECT  0.000 -0.330 0.270 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.570 2.070 2.000 2.730 ;
        RECT  1.460 1.735 1.570 2.730 ;
        RECT  0.445 2.070 1.460 2.730 ;
        RECT  0.335 1.800 0.445 2.730 ;
        RECT  0.000 2.070 0.335 2.730 ;
        END
    END VDD
END CELL108

MACRO CELL103
    CLASS CORE ;
    FOREIGN CELL103 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 2.400 ;
    SYMMETRY x y ;
    PIN ZN
        ANTENNADIFFAREA 0.2688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 0.510 3.350 1.890 ;
        RECT  3.225 0.510 3.250 0.890 ;
        RECT  3.225 1.310 3.250 1.890 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.1009 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.820 0.910 2.950 1.290 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1291 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.190 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 1.000 1.550 1.400 ;
        RECT  1.390 1.000 1.450 1.175 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.065 -0.330 3.400 0.330 ;
        RECT  2.955 -0.330 3.065 0.600 ;
        RECT  1.990 -0.330 2.955 0.330 ;
        RECT  1.890 -0.330 1.990 0.800 ;
        RECT  1.530 -0.330 1.890 0.330 ;
        RECT  1.420 -0.330 1.530 0.470 ;
        RECT  0.445 -0.330 1.420 0.330 ;
        RECT  0.335 -0.330 0.445 0.600 ;
        RECT  0.000 -0.330 0.335 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.055 2.070 3.400 2.730 ;
        RECT  2.945 1.800 3.055 2.730 ;
        RECT  2.045 2.070 2.945 2.730 ;
        RECT  1.955 1.435 2.045 2.730 ;
        RECT  1.850 1.435 1.955 1.545 ;
        RECT  0.470 2.070 1.955 2.730 ;
        RECT  0.360 1.600 0.470 2.730 ;
        RECT  0.000 2.070 0.360 2.730 ;
        END
    END VDD
END CELL103

MACRO CELL63
    CLASS CORE ;
    FOREIGN CELL63 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 0.2856 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 0.510 1.950 1.910 ;
        RECT  1.805 0.510 1.850 0.890 ;
        RECT  1.765 1.800 1.850 1.910 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.1009 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.710 1.560 1.160 ;
        RECT  1.375 0.990 1.450 1.160 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1311 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.995 0.375 1.400 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 -0.330 2.000 0.330 ;
        RECT  1.520 -0.330 1.630 0.600 ;
        RECT  0.365 -0.330 1.520 0.330 ;
        RECT  0.365 0.745 0.480 0.855 ;
        RECT  0.270 -0.330 0.365 0.855 ;
        RECT  0.000 -0.330 0.270 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 2.070 2.000 2.730 ;
        RECT  1.520 1.800 1.630 2.730 ;
        RECT  0.000 2.070 1.520 2.730 ;
        END
    END VDD
END CELL63

MACRO CELL11
    CLASS CORE ;
    FOREIGN CELL11 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.400 BY 2.400 ;
    SYMMETRY x y ;
    PIN Z
        ANTENNADIFFAREA 0.2688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 0.510 3.350 1.890 ;
        RECT  3.225 0.510 3.250 0.890 ;
        RECT  3.225 1.310 3.250 1.890 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.820 0.910 2.950 1.290 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.1024 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.050 0.910 0.190 1.290 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1008 ;
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 1.000 1.550 1.400 ;
        RECT  1.390 1.000 1.450 1.175 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.070 -0.330 3.400 0.330 ;
        RECT  2.960 -0.330 3.070 0.800 ;
        RECT  1.990 -0.330 2.960 0.330 ;
        RECT  1.890 -0.330 1.990 0.800 ;
        RECT  1.540 -0.330 1.890 0.330 ;
        RECT  1.430 -0.330 1.540 0.600 ;
        RECT  0.445 -0.330 1.430 0.330 ;
        RECT  0.335 -0.330 0.445 0.600 ;
        RECT  0.000 -0.330 0.335 0.330 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.045 2.070 3.400 2.730 ;
        RECT  2.935 1.800 3.045 2.730 ;
        RECT  2.045 2.070 2.935 2.730 ;
        RECT  1.955 1.435 2.045 2.730 ;
        RECT  1.850 1.435 1.955 1.545 ;
        RECT  0.470 2.070 1.955 2.730 ;
        RECT  0.360 1.600 0.470 2.730 ;
        RECT  0.000 2.070 0.360 2.730 ;
        END
    END VDD
END CELL11

END LIBRARY
